module layer_10_featuremap_213(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b83c725),
	.w1(32'h3ab06e20),
	.w2(32'h3c82116a),
	.w3(32'h3b1ca7ce),
	.w4(32'hbc5f4d52),
	.w5(32'h3b7374dd),
	.w6(32'h3c17f980),
	.w7(32'h3c162a68),
	.w8(32'hbb52ae64),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c16ae05),
	.w1(32'hbbe56744),
	.w2(32'hbc0135d8),
	.w3(32'h3c6dfea9),
	.w4(32'hbba4aa04),
	.w5(32'hbba860f3),
	.w6(32'hbc1c7b4e),
	.w7(32'hbbef3dc7),
	.w8(32'hbbcf768f),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7d5653),
	.w1(32'h3be3f5e7),
	.w2(32'hbb2528b4),
	.w3(32'hbb1740ba),
	.w4(32'h3a13ab21),
	.w5(32'hbb83065e),
	.w6(32'h3bbc490e),
	.w7(32'hb9e9ef22),
	.w8(32'hb9f6c15c),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1ff0f8),
	.w1(32'hbc9c4fac),
	.w2(32'hbbcadfb1),
	.w3(32'hba9662c4),
	.w4(32'h3aa93d57),
	.w5(32'hba54a14e),
	.w6(32'hbc85dbca),
	.w7(32'hbbea48bf),
	.w8(32'h3b9eb8f9),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b89feff),
	.w1(32'hbca9faa7),
	.w2(32'hbc00c25b),
	.w3(32'hbb13c4c3),
	.w4(32'hbc2a96e9),
	.w5(32'hbc410e77),
	.w6(32'hbc3820ae),
	.w7(32'hbc5b6fc7),
	.w8(32'h3c1c36b6),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9d8ac7),
	.w1(32'hbc48b9be),
	.w2(32'hbc2c5ac7),
	.w3(32'h3b3a5b34),
	.w4(32'hbc12f460),
	.w5(32'hbb9f8197),
	.w6(32'hbc3b4e41),
	.w7(32'hbc0073c8),
	.w8(32'hbac3ca71),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbec3d2a),
	.w1(32'hbc54bf34),
	.w2(32'hbcacf095),
	.w3(32'hbb2f3e88),
	.w4(32'hbc597660),
	.w5(32'hbcb46b9e),
	.w6(32'hbb54461d),
	.w7(32'hbc6ef6ec),
	.w8(32'hbc4bfc04),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc483cf),
	.w1(32'hbc1a75ea),
	.w2(32'hbb03e407),
	.w3(32'hbc9ce29f),
	.w4(32'hbbe8b45e),
	.w5(32'hbaac262d),
	.w6(32'hbc0ec762),
	.w7(32'hbb31604e),
	.w8(32'hba928f66),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb229cbd),
	.w1(32'hbab54b38),
	.w2(32'h3aebd349),
	.w3(32'h3a1ac21d),
	.w4(32'h399123f8),
	.w5(32'h3b921eda),
	.w6(32'hbafe26a6),
	.w7(32'h3b260fde),
	.w8(32'h3be4df95),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5aff0d),
	.w1(32'hbbf3b7e1),
	.w2(32'hbc4f4ab4),
	.w3(32'h3bc99461),
	.w4(32'hbb54005f),
	.w5(32'hbbd4a90e),
	.w6(32'hbb9f849a),
	.w7(32'hbaa39af5),
	.w8(32'hbbcae57b),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b6489),
	.w1(32'hbbb5fc5c),
	.w2(32'hbb7133ef),
	.w3(32'hbb7cae79),
	.w4(32'hba4249b4),
	.w5(32'h39c7c74e),
	.w6(32'hbc1b71c1),
	.w7(32'hbb1e8d8a),
	.w8(32'h3a9a7d7f),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba48901),
	.w1(32'hbbf622bd),
	.w2(32'hbc0ed784),
	.w3(32'hbc1f6db8),
	.w4(32'hba5b2d99),
	.w5(32'hbc49a7eb),
	.w6(32'hbc0b0e8c),
	.w7(32'hbb3fed1f),
	.w8(32'h3af2d577),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaff26d1),
	.w1(32'h3afa3b0e),
	.w2(32'hbb988a8c),
	.w3(32'hbc1951ca),
	.w4(32'h3bb18938),
	.w5(32'h39a90f5e),
	.w6(32'h3b11b3bf),
	.w7(32'h3bc0c7dc),
	.w8(32'h3ade7eae),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d28ca),
	.w1(32'h3b9fdaac),
	.w2(32'hbabdb5a6),
	.w3(32'hbaf157e8),
	.w4(32'h3b0b0e28),
	.w5(32'h3a492aea),
	.w6(32'h3c1171c9),
	.w7(32'h3b4c5aef),
	.w8(32'hbc094f44),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9f2a26),
	.w1(32'hbc7145ed),
	.w2(32'hbc2ca979),
	.w3(32'hbc328a72),
	.w4(32'h3c38d102),
	.w5(32'hbbc82838),
	.w6(32'hbcaa369a),
	.w7(32'hbc08a1be),
	.w8(32'h3c8fa570),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9170a6),
	.w1(32'hbbdf6ba7),
	.w2(32'hbc07abcc),
	.w3(32'hbc7df7f3),
	.w4(32'hba619ce9),
	.w5(32'h3ba155e4),
	.w6(32'hbc350888),
	.w7(32'hbaa4da8a),
	.w8(32'h3a5744ae),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbee31c),
	.w1(32'h3aa2481c),
	.w2(32'hbb2f0122),
	.w3(32'h3bbef8d8),
	.w4(32'hbb6b28d5),
	.w5(32'hba1fa945),
	.w6(32'hbb5037f8),
	.w7(32'hbb22c99b),
	.w8(32'hb84de8bb),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc074c4f),
	.w1(32'hbbef3459),
	.w2(32'hbc1a5710),
	.w3(32'h391daa9a),
	.w4(32'hbb2870e6),
	.w5(32'hbb7e0990),
	.w6(32'hbc066871),
	.w7(32'h3a6a538e),
	.w8(32'h3ba73201),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9890b3),
	.w1(32'h3ab1f1ea),
	.w2(32'hbb7e9c9f),
	.w3(32'h3afb28e6),
	.w4(32'h3b4eab2e),
	.w5(32'hbb3827c1),
	.w6(32'h38f8d86f),
	.w7(32'h3b649ca0),
	.w8(32'h3b099a88),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a64c4d3),
	.w1(32'hba6fa6e3),
	.w2(32'hbad4650f),
	.w3(32'hb9b74cd8),
	.w4(32'hba5b3f34),
	.w5(32'h3ac33ed8),
	.w6(32'hbae21871),
	.w7(32'hba0f6850),
	.w8(32'h3b4de899),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8e5d25),
	.w1(32'hbb493f8d),
	.w2(32'hbbe600bf),
	.w3(32'h3b9d95c8),
	.w4(32'hba246ace),
	.w5(32'hb89f0af1),
	.w6(32'hbb2da90f),
	.w7(32'hbb1df2ed),
	.w8(32'h38e2e88a),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7daf4d),
	.w1(32'h3c13413b),
	.w2(32'hb942763e),
	.w3(32'h3a97a190),
	.w4(32'hbc7091fb),
	.w5(32'hbb9a45ca),
	.w6(32'h3b5ac8e0),
	.w7(32'h3b64e461),
	.w8(32'hbc2393fa),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5c908a),
	.w1(32'hbbf8a22b),
	.w2(32'hbc5a6d13),
	.w3(32'h3a109870),
	.w4(32'hbb4b6e28),
	.w5(32'hbbfdb52b),
	.w6(32'hbc386ae4),
	.w7(32'hbc022768),
	.w8(32'hbc60a9b1),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4f88a6),
	.w1(32'hbb003e73),
	.w2(32'hbc01bc8d),
	.w3(32'h3c117d29),
	.w4(32'h3856e5fa),
	.w5(32'hbb73e556),
	.w6(32'hbaa07667),
	.w7(32'h3aeb81b7),
	.w8(32'hbb5b635e),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb33f2ef),
	.w1(32'hbc4c197a),
	.w2(32'hbb40b60c),
	.w3(32'hbb1ed6f1),
	.w4(32'hbab38e2e),
	.w5(32'h3a10177b),
	.w6(32'hbc66a2a3),
	.w7(32'hba02f28c),
	.w8(32'hba82fbdc),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba9dc20),
	.w1(32'h3b98f198),
	.w2(32'hba8c395b),
	.w3(32'h3af11f42),
	.w4(32'hbc6516de),
	.w5(32'hbbd0e0b9),
	.w6(32'h3b8a2ec4),
	.w7(32'hbabfad93),
	.w8(32'hbc562a5c),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe30431),
	.w1(32'h3ab4e4ea),
	.w2(32'hbb0ada07),
	.w3(32'h39f61695),
	.w4(32'hba2f80bb),
	.w5(32'h3aa29c92),
	.w6(32'h3a0d7da1),
	.w7(32'hba5819be),
	.w8(32'h3afa6f9c),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b74c031),
	.w1(32'hbb054924),
	.w2(32'h3b8607a6),
	.w3(32'h3b0b475d),
	.w4(32'h3bc43e8f),
	.w5(32'h3baeb211),
	.w6(32'hbb2eb52b),
	.w7(32'h3c19586a),
	.w8(32'h3bcc4b52),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b95c757),
	.w1(32'h3ba359ae),
	.w2(32'hbad91bff),
	.w3(32'hbb1b882d),
	.w4(32'h3bc28c89),
	.w5(32'hbaaf1808),
	.w6(32'h3c1335fc),
	.w7(32'h3b75eada),
	.w8(32'h3ba86fb6),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcef0e9),
	.w1(32'h3bb8adbd),
	.w2(32'h3b37c694),
	.w3(32'h3ae7ccf5),
	.w4(32'h39be488f),
	.w5(32'hbb211a03),
	.w6(32'hb9e7e6fc),
	.w7(32'h3b010503),
	.w8(32'hba40833e),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb12552),
	.w1(32'hbacc6f6c),
	.w2(32'hbb71e438),
	.w3(32'h39d20f70),
	.w4(32'hb9da1f8a),
	.w5(32'hb9dd2db2),
	.w6(32'hbae1d413),
	.w7(32'hbb077d63),
	.w8(32'h3992e791),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37c9eee7),
	.w1(32'h3a59b981),
	.w2(32'hbab5ff3e),
	.w3(32'h3aa7b821),
	.w4(32'hb9af44b9),
	.w5(32'h3a6ae18c),
	.w6(32'h3a00fbad),
	.w7(32'hba66dbc6),
	.w8(32'h3a46210f),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0bda1b),
	.w1(32'hbba5fb83),
	.w2(32'hbd039100),
	.w3(32'h3aced0a7),
	.w4(32'hbbbd73e8),
	.w5(32'hbcf7b0fe),
	.w6(32'hbbaa78e3),
	.w7(32'hbd0208ec),
	.w8(32'hbc956d35),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb10dee),
	.w1(32'h3d29bdd7),
	.w2(32'h3ca2a10f),
	.w3(32'hbca3dbdc),
	.w4(32'h3c46739c),
	.w5(32'h3c43eb02),
	.w6(32'h3cb4fe4e),
	.w7(32'h3b3691b1),
	.w8(32'hbafe9cd2),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1d0ae8),
	.w1(32'hbb54ff6e),
	.w2(32'h3b93c152),
	.w3(32'h3bb360d5),
	.w4(32'hbb72fda7),
	.w5(32'h3ba18f5d),
	.w6(32'hbb7fdbfe),
	.w7(32'h3bd574cd),
	.w8(32'h3c37cb40),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2aef5f),
	.w1(32'hbbd0cd0d),
	.w2(32'hbbc02a09),
	.w3(32'h3c0943d0),
	.w4(32'hbb1a6edb),
	.w5(32'hba374d6f),
	.w6(32'hbaf865bf),
	.w7(32'hbb3b26a0),
	.w8(32'hba8b6162),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc822299),
	.w1(32'hbcbdac34),
	.w2(32'hbc709ee9),
	.w3(32'hbbed78a8),
	.w4(32'hbc4768c4),
	.w5(32'hbc28b938),
	.w6(32'hbc3b4f83),
	.w7(32'hbc1bf30f),
	.w8(32'hbb9e328b),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6eba5a),
	.w1(32'h3b39bef1),
	.w2(32'hbbe5d865),
	.w3(32'hbbe9f10a),
	.w4(32'h3a490728),
	.w5(32'hbbae83cb),
	.w6(32'hbc2d0c5a),
	.w7(32'hbc167033),
	.w8(32'hbc34a4f4),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1e539f),
	.w1(32'hba34019c),
	.w2(32'hbbcc7427),
	.w3(32'hbbc440f7),
	.w4(32'hbbe42192),
	.w5(32'hbc110a92),
	.w6(32'hbbb530aa),
	.w7(32'hbbcc9aae),
	.w8(32'hbc2526ad),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b57ba97),
	.w1(32'hbb08cddb),
	.w2(32'hbb7f90ef),
	.w3(32'h3b6a75bd),
	.w4(32'hba2eb577),
	.w5(32'hbb315534),
	.w6(32'hbb8e55d2),
	.w7(32'hbb536d57),
	.w8(32'hb905afde),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cee5f8),
	.w1(32'h3ba0aee7),
	.w2(32'h3bd09a16),
	.w3(32'hba326182),
	.w4(32'h3b7063fd),
	.w5(32'h3b0054b1),
	.w6(32'h3bbbc307),
	.w7(32'h3ba38e8a),
	.w8(32'h3bac501a),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf96501),
	.w1(32'hb8caf849),
	.w2(32'h3a7e1801),
	.w3(32'h3b1771fb),
	.w4(32'h3b88a41b),
	.w5(32'h3b364ca3),
	.w6(32'hbb495ab4),
	.w7(32'hbb437c84),
	.w8(32'h3b58f26a),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b24e358),
	.w1(32'h3b8bc79e),
	.w2(32'hba74df20),
	.w3(32'hbba12bbe),
	.w4(32'h39cb63a1),
	.w5(32'hbaa64e7c),
	.w6(32'hbb205d7f),
	.w7(32'hbb2ec0f0),
	.w8(32'hba8d2693),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc02cf32),
	.w1(32'hbc0fd596),
	.w2(32'hbb95e217),
	.w3(32'hbb892826),
	.w4(32'hbb01b359),
	.w5(32'hba1a613f),
	.w6(32'hbbfe1165),
	.w7(32'h3bf2a424),
	.w8(32'hbb5dc741),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb857905),
	.w1(32'h3c6c1b1f),
	.w2(32'h3afe9fd5),
	.w3(32'hbb27a5bb),
	.w4(32'h3c15155e),
	.w5(32'h3bcbc26e),
	.w6(32'h3c1f5183),
	.w7(32'h3bbba53d),
	.w8(32'hbc5cce92),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8c6163),
	.w1(32'hbb5f2c49),
	.w2(32'hbc72bdbf),
	.w3(32'h3b261f52),
	.w4(32'h39bf5faf),
	.w5(32'hbbbc03ca),
	.w6(32'hbb96e383),
	.w7(32'hbc11513e),
	.w8(32'hbc5a9ab6),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc207687),
	.w1(32'hbbba79e7),
	.w2(32'hbc2dc25a),
	.w3(32'hbb1cfbeb),
	.w4(32'h3bbd4350),
	.w5(32'hbb8bf561),
	.w6(32'hbc37f046),
	.w7(32'hbbef5597),
	.w8(32'h3b9ab449),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3999dc9c),
	.w1(32'h3b9b751e),
	.w2(32'h3a72a3bc),
	.w3(32'hbbf36f18),
	.w4(32'h3b9b7b0b),
	.w5(32'h3bddaf6b),
	.w6(32'h3bec5901),
	.w7(32'h3c7dfe04),
	.w8(32'h3c43af82),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1a8912),
	.w1(32'h3b72f953),
	.w2(32'hba719a21),
	.w3(32'h3c2968bb),
	.w4(32'h3934298a),
	.w5(32'hb9e1fc1e),
	.w6(32'h3a7c3cd0),
	.w7(32'hbb0fe7ce),
	.w8(32'h3ad00bf7),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c3c9b1),
	.w1(32'hbae99fc5),
	.w2(32'hbb46c588),
	.w3(32'h3a4eb9ff),
	.w4(32'hbb31533d),
	.w5(32'hbb2798ea),
	.w6(32'hb89245c9),
	.w7(32'hba2dde3d),
	.w8(32'hbb2e9231),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c5145),
	.w1(32'h3bf55744),
	.w2(32'hbbb4372e),
	.w3(32'hbadf51fc),
	.w4(32'h3bbcb8d2),
	.w5(32'hbb977fa0),
	.w6(32'h3c0e50e8),
	.w7(32'h3ab7338b),
	.w8(32'hbbd282dd),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc83290a),
	.w1(32'hbc0055b6),
	.w2(32'h3c72d869),
	.w3(32'hbc31d0bb),
	.w4(32'h3bd03413),
	.w5(32'h3c2b6c6d),
	.w6(32'hbc13a844),
	.w7(32'h3bba44e4),
	.w8(32'h3c63ad24),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3c9a15),
	.w1(32'hbba4d54e),
	.w2(32'hbc5bf042),
	.w3(32'hb6fc7b8e),
	.w4(32'hbb2728d3),
	.w5(32'hbb287a19),
	.w6(32'hbbac2849),
	.w7(32'hbba79ce4),
	.w8(32'h3aa4c70b),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc23c80a),
	.w1(32'hbcda91bb),
	.w2(32'hbc97a9e6),
	.w3(32'hba0ea732),
	.w4(32'hbc7d707a),
	.w5(32'hbc8d42c5),
	.w6(32'hbc88cc22),
	.w7(32'hbc2422e0),
	.w8(32'hbb30339b),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabb20a1),
	.w1(32'hbac73f84),
	.w2(32'hbb62a6d6),
	.w3(32'h3b820329),
	.w4(32'h386c3590),
	.w5(32'hbb0c2c81),
	.w6(32'hb9851e68),
	.w7(32'hb9706055),
	.w8(32'hbaf02a7f),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaebd51e),
	.w1(32'hbbc7733e),
	.w2(32'hbbdc63fa),
	.w3(32'hb9be190f),
	.w4(32'h3ade3a35),
	.w5(32'hbc21d9a0),
	.w6(32'hbb1c59b1),
	.w7(32'hbb891865),
	.w8(32'hbae3e98a),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3e698d),
	.w1(32'h3c29174c),
	.w2(32'hbba9caa8),
	.w3(32'hbbc9925d),
	.w4(32'h3c60ef96),
	.w5(32'h3abbd280),
	.w6(32'h3bda6472),
	.w7(32'h3a25e4cf),
	.w8(32'hbac4ce70),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc37b76),
	.w1(32'hbc941bc0),
	.w2(32'hbb8472a5),
	.w3(32'hbb3bf0d5),
	.w4(32'hbc158164),
	.w5(32'hbc61543e),
	.w6(32'hbbe51f62),
	.w7(32'hbc5697be),
	.w8(32'hbbca096f),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc88d86d),
	.w1(32'hb99af234),
	.w2(32'h3b57487f),
	.w3(32'hbc252133),
	.w4(32'hba5f3931),
	.w5(32'h3b0a90f7),
	.w6(32'h397a7ccb),
	.w7(32'h3ba4550e),
	.w8(32'h3b6700a3),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba4c80b),
	.w1(32'h3947fd47),
	.w2(32'h3862e825),
	.w3(32'h3b464f19),
	.w4(32'hbb58646a),
	.w5(32'h3a083292),
	.w6(32'hb9427f3d),
	.w7(32'h3a3f455b),
	.w8(32'h3ad67758),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7d7292),
	.w1(32'hbaca8498),
	.w2(32'hbb35bea2),
	.w3(32'h3adca72d),
	.w4(32'hba5eb334),
	.w5(32'hbb2338a7),
	.w6(32'hba3a83ff),
	.w7(32'h3b60d242),
	.w8(32'hbae3a7ef),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdf61f4),
	.w1(32'h3b0d6b6d),
	.w2(32'hbb78a045),
	.w3(32'hbb5de6ed),
	.w4(32'hba9f6112),
	.w5(32'h39d666ee),
	.w6(32'h3a98cabe),
	.w7(32'h3b7b5358),
	.w8(32'hbb1b8bfc),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2f8458),
	.w1(32'hbb67606f),
	.w2(32'hbc6b6613),
	.w3(32'h3b654ee4),
	.w4(32'hbc1cad69),
	.w5(32'hbcca26c9),
	.w6(32'hbb8d96c4),
	.w7(32'hbcb7e81a),
	.w8(32'hbbc2066d),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdfd183),
	.w1(32'hbbb3afe4),
	.w2(32'h3b127566),
	.w3(32'hbb479876),
	.w4(32'hbb739bf3),
	.w5(32'h3a98090e),
	.w6(32'hbb950c62),
	.w7(32'h3af3f220),
	.w8(32'h39f09361),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8832b4d),
	.w1(32'h3a6884a0),
	.w2(32'hbb8faeb5),
	.w3(32'hba9f9b8a),
	.w4(32'h3b1eaa4b),
	.w5(32'hbb65d95f),
	.w6(32'h3a00fc00),
	.w7(32'hbbb95508),
	.w8(32'hbb0e5937),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ce3a9),
	.w1(32'h3b37bb4b),
	.w2(32'h3c08f50c),
	.w3(32'hbbd62964),
	.w4(32'h3b67b94c),
	.w5(32'hba539714),
	.w6(32'h3acf8da5),
	.w7(32'hbb3d8d48),
	.w8(32'hbc00d07c),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9cd925),
	.w1(32'h3b63dfc8),
	.w2(32'hbb0c2409),
	.w3(32'hbc6c9af2),
	.w4(32'hb48dacb0),
	.w5(32'hbb3b7ae0),
	.w6(32'hbb4f604d),
	.w7(32'h3b0e287f),
	.w8(32'hba902310),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3a19fc),
	.w1(32'hbc14ccde),
	.w2(32'hbc3c94ca),
	.w3(32'hbbcfcdb7),
	.w4(32'hbb1dccbf),
	.w5(32'hbc10a123),
	.w6(32'hba8bfe7a),
	.w7(32'hbbcd369b),
	.w8(32'hbb89db24),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe59a95),
	.w1(32'hbbbda787),
	.w2(32'hbc415225),
	.w3(32'h3b032354),
	.w4(32'hba1a8db8),
	.w5(32'hbac93c47),
	.w6(32'hbbf79aba),
	.w7(32'hbafe9c5f),
	.w8(32'hba632b68),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be6e6d5),
	.w1(32'h3a8897b3),
	.w2(32'hbcc3a41b),
	.w3(32'h3b9bcf35),
	.w4(32'h3c206793),
	.w5(32'hbc8a9bc4),
	.w6(32'hbbbaff12),
	.w7(32'hbc11e06a),
	.w8(32'hbce193f8),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce0cce9),
	.w1(32'hbaa3caae),
	.w2(32'h3b4d8dbf),
	.w3(32'hbc978b3f),
	.w4(32'h3a1da498),
	.w5(32'h3b431fab),
	.w6(32'hbada4709),
	.w7(32'h3bb25685),
	.w8(32'h3c1daffa),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2a8135),
	.w1(32'hbb931356),
	.w2(32'h3a430f86),
	.w3(32'h3b95a715),
	.w4(32'hbb3e8b6e),
	.w5(32'h3b0e49ef),
	.w6(32'hbb61bf79),
	.w7(32'h3aa01076),
	.w8(32'h3b879fb5),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b96305a),
	.w1(32'hbb029b9d),
	.w2(32'hb9bb2e42),
	.w3(32'h3b7023b9),
	.w4(32'hbb14a802),
	.w5(32'h3a645e4d),
	.w6(32'hba9adfff),
	.w7(32'h3ad03b79),
	.w8(32'h3b5cbf4a),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b11e20b),
	.w1(32'hbaf651f2),
	.w2(32'hbb8df09d),
	.w3(32'h3b1fd059),
	.w4(32'hba83cfe4),
	.w5(32'h3aaefb70),
	.w6(32'hbac690ff),
	.w7(32'hbaad883d),
	.w8(32'h398b12fc),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa37d6a),
	.w1(32'hbbbcc715),
	.w2(32'h3a435c7f),
	.w3(32'h3ade6986),
	.w4(32'hb8b25a26),
	.w5(32'h39fb7d0c),
	.w6(32'hbbc275da),
	.w7(32'hba614a57),
	.w8(32'h3b30416f),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8135e8),
	.w1(32'hbaf027a1),
	.w2(32'hbba5e68a),
	.w3(32'hbbac222d),
	.w4(32'h3b9065f6),
	.w5(32'hbc1c36e1),
	.w6(32'hbc0aa1b0),
	.w7(32'hbbc860df),
	.w8(32'h3af65b6d),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4d3162),
	.w1(32'hbbd490fc),
	.w2(32'hbb958103),
	.w3(32'hbca2b880),
	.w4(32'hbbb9cb61),
	.w5(32'h3acd2c39),
	.w6(32'hbb525878),
	.w7(32'hba08b2d4),
	.w8(32'hbb6e2d91),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1fc4fe),
	.w1(32'h3b6ef3e8),
	.w2(32'h3c42e0f9),
	.w3(32'hbb0fed2b),
	.w4(32'h3bdb7354),
	.w5(32'h3be59d30),
	.w6(32'h3b180a3b),
	.w7(32'h3c39148f),
	.w8(32'hb9f947e9),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad8e1e1),
	.w1(32'hbba67b76),
	.w2(32'hbb52ff33),
	.w3(32'h3ae9a99c),
	.w4(32'hbb5a3262),
	.w5(32'hbb3ef959),
	.w6(32'hbb182450),
	.w7(32'hbb295cb7),
	.w8(32'hbba97b6b),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbda9c39),
	.w1(32'hbad6c8d9),
	.w2(32'hbbeba649),
	.w3(32'h3ab65925),
	.w4(32'hbaba729a),
	.w5(32'hbb2199a9),
	.w6(32'hbaf13e31),
	.w7(32'hba93ef8c),
	.w8(32'h3a9db208),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38303ef5),
	.w1(32'hbb0c4c29),
	.w2(32'hbc31f9e6),
	.w3(32'h3acfb522),
	.w4(32'h3b00df31),
	.w5(32'hbbb78aac),
	.w6(32'h3b2b8b47),
	.w7(32'hba622665),
	.w8(32'hb9a319b5),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb233f35),
	.w1(32'h3bf8bbe0),
	.w2(32'hbc08cac9),
	.w3(32'h3a9975de),
	.w4(32'h3bb48ff5),
	.w5(32'hbaa47e10),
	.w6(32'h3b9331ef),
	.w7(32'hbaa9edad),
	.w8(32'hbb3a5d8f),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc338b2),
	.w1(32'hbbd1237e),
	.w2(32'hba1e1665),
	.w3(32'hbac0da9f),
	.w4(32'hbb28d67c),
	.w5(32'h3a8d843e),
	.w6(32'hbb4e9b56),
	.w7(32'h3b4bff6c),
	.w8(32'h3c0ce99f),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c066240),
	.w1(32'hba24b676),
	.w2(32'h3acd0a3c),
	.w3(32'h3b948041),
	.w4(32'hbb31c3e5),
	.w5(32'h38594414),
	.w6(32'h3b27e138),
	.w7(32'h3b1d5f57),
	.w8(32'hbb0be3e7),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3937b14f),
	.w1(32'h3b1a3d81),
	.w2(32'h3a0f69d6),
	.w3(32'h39d74dc3),
	.w4(32'h3a887d82),
	.w5(32'hb7d768bd),
	.w6(32'hb9993f15),
	.w7(32'h3a5700af),
	.w8(32'hbb229ee8),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a888253),
	.w1(32'h3b5aaa2c),
	.w2(32'hbb968249),
	.w3(32'hba9ba1d5),
	.w4(32'h3b5d4a17),
	.w5(32'hbac1da91),
	.w6(32'h3b2e8d2f),
	.w7(32'hbb3f45d9),
	.w8(32'hbb2af46d),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc2144c),
	.w1(32'h3bfcc617),
	.w2(32'h3c913fb3),
	.w3(32'hbb7c77f9),
	.w4(32'h3c20ff59),
	.w5(32'h3c45140a),
	.w6(32'h3bc7d0cf),
	.w7(32'h3c8b4e81),
	.w8(32'hbb268b43),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8e865b),
	.w1(32'hba4a544f),
	.w2(32'hbb5675fa),
	.w3(32'h39ae27dc),
	.w4(32'hb52673d2),
	.w5(32'h3a6820fa),
	.w6(32'hbaf0697f),
	.w7(32'hbabd782d),
	.w8(32'h3a5026fa),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb05c99a),
	.w1(32'hbb3a3859),
	.w2(32'hbbb47395),
	.w3(32'h3ac2d59d),
	.w4(32'h39bd11a9),
	.w5(32'hbb76e5e4),
	.w6(32'hbb57fba0),
	.w7(32'hbadf5fc6),
	.w8(32'hbb70b713),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5d87ee),
	.w1(32'hbbbb4cc8),
	.w2(32'hbc0e2409),
	.w3(32'hbc230d9c),
	.w4(32'hb9e3b4fb),
	.w5(32'hbb1fcd12),
	.w6(32'hbc3ac3c4),
	.w7(32'hbbb1e180),
	.w8(32'hba7b53fa),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b88c4cc),
	.w1(32'h3a3148fc),
	.w2(32'hbb9b148c),
	.w3(32'h3b278b3c),
	.w4(32'hbb3ffd08),
	.w5(32'hbba1801f),
	.w6(32'hbaa85329),
	.w7(32'hbaae3b44),
	.w8(32'hbb40fae2),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd7aaba),
	.w1(32'hbb27fc70),
	.w2(32'hbc3ada65),
	.w3(32'hbb8c4205),
	.w4(32'hbb5b1c80),
	.w5(32'hbc1d8042),
	.w6(32'hbb4e217c),
	.w7(32'hbc254341),
	.w8(32'hbc50b418),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1a450a),
	.w1(32'hbb4dafaa),
	.w2(32'hbc02c22b),
	.w3(32'hbbdfddca),
	.w4(32'hbba120f4),
	.w5(32'hbbf03903),
	.w6(32'hbb8edf54),
	.w7(32'h3ae7b7d8),
	.w8(32'h3b1af053),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe7e653),
	.w1(32'hbbb99058),
	.w2(32'hbc62abd8),
	.w3(32'hbbc0b087),
	.w4(32'h3b5bc5ca),
	.w5(32'hbb0c81a6),
	.w6(32'hbb5d0f78),
	.w7(32'hbb8b5ad4),
	.w8(32'h3a70fa0f),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba99522b),
	.w1(32'hba1c5df4),
	.w2(32'hbb9842b8),
	.w3(32'h39d339ec),
	.w4(32'hbb8c44e3),
	.w5(32'hbba7497c),
	.w6(32'hb9c298d6),
	.w7(32'h39b96cf0),
	.w8(32'hbb915eb8),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adecb99),
	.w1(32'hbc107e5e),
	.w2(32'hbc2cd75e),
	.w3(32'hb99b57d1),
	.w4(32'hbc718824),
	.w5(32'hbc43c9d5),
	.w6(32'hbbd8f56c),
	.w7(32'hbc0264f1),
	.w8(32'hbc02764d),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2368eb),
	.w1(32'h3999b1a2),
	.w2(32'h3a86d2ec),
	.w3(32'h3b5a80c2),
	.w4(32'hbb291eb0),
	.w5(32'hbb1cf069),
	.w6(32'h3b32b110),
	.w7(32'hba7d32bd),
	.w8(32'h3b14629b),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b7d3af),
	.w1(32'hbc009b28),
	.w2(32'hbbdfd018),
	.w3(32'h3b3e8120),
	.w4(32'hbb2ea351),
	.w5(32'hbba864e3),
	.w6(32'hbbffa6ce),
	.w7(32'hbbc855b0),
	.w8(32'hbb829dd1),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390ba08a),
	.w1(32'h3b45e88b),
	.w2(32'hbc2ba1c6),
	.w3(32'h3b07b31a),
	.w4(32'hba44dd58),
	.w5(32'hbbf98da1),
	.w6(32'h3ba5c75f),
	.w7(32'hba06fa64),
	.w8(32'hb9474c59),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcafe978),
	.w1(32'hbc9a6a9f),
	.w2(32'hbc228e69),
	.w3(32'hbc0ad683),
	.w4(32'hbbb95dfa),
	.w5(32'h3b134c4f),
	.w6(32'hbbecabe3),
	.w7(32'h3a7d5b3e),
	.w8(32'h39dbc204),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5cb887),
	.w1(32'hbb64e099),
	.w2(32'hbaea4e25),
	.w3(32'h3a2673c9),
	.w4(32'h3b512f05),
	.w5(32'hbbc74a59),
	.w6(32'hbb17668c),
	.w7(32'hbc833058),
	.w8(32'hbbc0ca9f),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3fde23),
	.w1(32'hbbe83b38),
	.w2(32'hbbffd8e2),
	.w3(32'hbbd968cd),
	.w4(32'hbc2e10f0),
	.w5(32'hbc496388),
	.w6(32'hbb4a47bb),
	.w7(32'hbc8149eb),
	.w8(32'hbc1d8f65),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1e4bc4),
	.w1(32'hbbc67b0d),
	.w2(32'hbbd3cece),
	.w3(32'h3c51c418),
	.w4(32'hbc0f2ad7),
	.w5(32'hbb85173c),
	.w6(32'h3b72cb08),
	.w7(32'hba07fb27),
	.w8(32'hbc212863),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc366a1c),
	.w1(32'hbbc8872d),
	.w2(32'hbb49c382),
	.w3(32'hbb2b25a0),
	.w4(32'hbb6d942b),
	.w5(32'h388dacfa),
	.w6(32'hbb8f7691),
	.w7(32'hba15fb9d),
	.w8(32'h3b8ebcea),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8b59c5),
	.w1(32'hbc60e412),
	.w2(32'hbc330108),
	.w3(32'hbbe3864e),
	.w4(32'hbc06f823),
	.w5(32'hbbab219d),
	.w6(32'hbbbd9d0c),
	.w7(32'h3b11bb1d),
	.w8(32'hbabdec06),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc010c1f),
	.w1(32'hbbc38709),
	.w2(32'hbc0e1b70),
	.w3(32'hbafe2616),
	.w4(32'hbba81310),
	.w5(32'hbbc56453),
	.w6(32'h38bea06e),
	.w7(32'hbb8041e1),
	.w8(32'hbb03dfdf),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a432428),
	.w1(32'h3c15860a),
	.w2(32'h3aeb5025),
	.w3(32'h3b2770dc),
	.w4(32'h3b7e10e7),
	.w5(32'h3a6468cf),
	.w6(32'h3c06a403),
	.w7(32'h3b901d2b),
	.w8(32'hb9e807eb),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e2314),
	.w1(32'hbbc71860),
	.w2(32'hbc1ee747),
	.w3(32'hbbdbfdfe),
	.w4(32'hbb933865),
	.w5(32'hbb06840a),
	.w6(32'hbb8ed42c),
	.w7(32'hbb996735),
	.w8(32'hbb552b18),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb558733),
	.w1(32'hb84d13d2),
	.w2(32'hbb7073be),
	.w3(32'h3b280fb8),
	.w4(32'hb8db17d9),
	.w5(32'hb9ea2fd8),
	.w6(32'h39b63495),
	.w7(32'h39a273fa),
	.w8(32'hbbc852d4),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb3f7b4),
	.w1(32'h3c3da56b),
	.w2(32'h3c02132d),
	.w3(32'hbaaf02b0),
	.w4(32'h3c224755),
	.w5(32'h3b602d63),
	.w6(32'h3bf2253b),
	.w7(32'h3b8a5ae6),
	.w8(32'hbbaba3eb),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc060b4a),
	.w1(32'hbb1b36d7),
	.w2(32'hbb6fadc8),
	.w3(32'hbb1b70af),
	.w4(32'hba0a624f),
	.w5(32'h3ac1d53c),
	.w6(32'hbb13c433),
	.w7(32'h39d4fcc7),
	.w8(32'h3ae20f36),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc8cf92),
	.w1(32'h3c14d236),
	.w2(32'h3d146ba3),
	.w3(32'h3bc8a876),
	.w4(32'h3beba8a8),
	.w5(32'h3cb2014d),
	.w6(32'h3be37b69),
	.w7(32'h3c5b747c),
	.w8(32'h3bd3bd77),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c46a7f1),
	.w1(32'hbbf905e7),
	.w2(32'hbb1a5733),
	.w3(32'h3c76efe6),
	.w4(32'h3a68ae79),
	.w5(32'h3b98cc71),
	.w6(32'hbc12893e),
	.w7(32'hbac38f0f),
	.w8(32'h3b82625e),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba605d5b),
	.w1(32'hbaa9476e),
	.w2(32'h3a8087e2),
	.w3(32'hbaad693e),
	.w4(32'h3b7de6df),
	.w5(32'h3bb0e9cc),
	.w6(32'hbba81e35),
	.w7(32'h3aebe810),
	.w8(32'h3a3a36a1),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b986d1c),
	.w1(32'h3c213755),
	.w2(32'h3b1522ff),
	.w3(32'hba4ee4c1),
	.w4(32'h3c406967),
	.w5(32'h3bd822de),
	.w6(32'h3bca2b0b),
	.w7(32'h3b96c7f3),
	.w8(32'hba9c7ca1),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdb678c),
	.w1(32'hbb204816),
	.w2(32'hbb382c2c),
	.w3(32'h39533780),
	.w4(32'hbb978a19),
	.w5(32'hbac619fb),
	.w6(32'h3a681f05),
	.w7(32'hb9d88577),
	.w8(32'hbb9e56eb),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1c9d60),
	.w1(32'hbb16157c),
	.w2(32'hbaa30e21),
	.w3(32'hbb483cf0),
	.w4(32'hbaf8ecb5),
	.w5(32'hbaa66c2e),
	.w6(32'hbb536323),
	.w7(32'hba89a73d),
	.w8(32'hba0169d9),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad3b7c4),
	.w1(32'hbb9ef05f),
	.w2(32'hbaef72ce),
	.w3(32'hba25c445),
	.w4(32'hbb85de18),
	.w5(32'hba853520),
	.w6(32'hbb851b28),
	.w7(32'hba294c2f),
	.w8(32'h3a94834f),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb85ae9e5),
	.w1(32'h3c2244e2),
	.w2(32'hb9f3a14f),
	.w3(32'h39f00ad2),
	.w4(32'hbbbc6d01),
	.w5(32'h3b79e729),
	.w6(32'h3be734b7),
	.w7(32'hbb066910),
	.w8(32'hbc376bff),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc298289),
	.w1(32'hbb16d795),
	.w2(32'hbb9e0e93),
	.w3(32'h3baebd9a),
	.w4(32'h3b16a0db),
	.w5(32'hbb712ed6),
	.w6(32'hbb3f349f),
	.w7(32'hbb058954),
	.w8(32'hbb7d2ff4),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb903b90),
	.w1(32'hbb853510),
	.w2(32'hbbb63dc9),
	.w3(32'hbaec9404),
	.w4(32'hba3a9502),
	.w5(32'hbabce259),
	.w6(32'hbb7939a6),
	.w7(32'hbb50def5),
	.w8(32'h3aa0bb64),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab13063),
	.w1(32'hbbc0f251),
	.w2(32'h39bf36d6),
	.w3(32'h3b513b06),
	.w4(32'hbb51c742),
	.w5(32'h3b86aace),
	.w6(32'hbafbd924),
	.w7(32'h3c046f73),
	.w8(32'h3bea5468),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0a9ee6),
	.w1(32'hbaee1367),
	.w2(32'hba3f48cc),
	.w3(32'h3ba818b0),
	.w4(32'hbb902c6f),
	.w5(32'hbb1a2b16),
	.w6(32'hbbfa9a8c),
	.w7(32'hbc0067c6),
	.w8(32'hbc15bb99),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4a0b0a),
	.w1(32'h3baa37fa),
	.w2(32'hbb01ba0e),
	.w3(32'h3a6c85da),
	.w4(32'hbc712e0b),
	.w5(32'h3b27cf24),
	.w6(32'h3c20e7e1),
	.w7(32'hbbe5eba9),
	.w8(32'hbc6936b4),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb48a834),
	.w1(32'hbc09ba77),
	.w2(32'hbc453aeb),
	.w3(32'h3c3d7719),
	.w4(32'hbbeb445d),
	.w5(32'hbbd51791),
	.w6(32'hbbe9536f),
	.w7(32'hbb18a0b4),
	.w8(32'h3b7fb769),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb25d3b2),
	.w1(32'hbb930f9f),
	.w2(32'hbb1a62bb),
	.w3(32'h39ea7e85),
	.w4(32'hbb29895a),
	.w5(32'h3b2a2d2a),
	.w6(32'hbb3a1091),
	.w7(32'h3a9ce600),
	.w8(32'h3b321226),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a92a5c2),
	.w1(32'h3a9b50de),
	.w2(32'h3a464272),
	.w3(32'h3b61b7e2),
	.w4(32'h3ab0030d),
	.w5(32'h3ac3f075),
	.w6(32'hba010ee8),
	.w7(32'hbac5624c),
	.w8(32'hbaad3810),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbab79c0),
	.w1(32'hbc14483a),
	.w2(32'hbbd9c053),
	.w3(32'h3a27dbef),
	.w4(32'hbb5bff34),
	.w5(32'hba1174ca),
	.w6(32'h3aaa1c0c),
	.w7(32'hbc01e287),
	.w8(32'hbba9c61a),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0a9c6b),
	.w1(32'hbc344695),
	.w2(32'hbc93cfa6),
	.w3(32'h3addbb55),
	.w4(32'hbb72dcd8),
	.w5(32'hbc1b3fb2),
	.w6(32'hbc3ae77c),
	.w7(32'hbc125cf4),
	.w8(32'hbc3513b3),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6389d3),
	.w1(32'hbc0b61a2),
	.w2(32'hbbd2751d),
	.w3(32'hbc38df14),
	.w4(32'hbbee9707),
	.w5(32'hbba1e72e),
	.w6(32'hbbff99d2),
	.w7(32'hbbde5135),
	.w8(32'hbbd5eecc),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2a4238),
	.w1(32'hbbe10713),
	.w2(32'hbb6c4df0),
	.w3(32'hbbdaaaf8),
	.w4(32'hbb096d19),
	.w5(32'hb9ec1e7a),
	.w6(32'hbbc9d0ed),
	.w7(32'hbba6993b),
	.w8(32'hbb3340ca),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb35f498),
	.w1(32'hbbfb5e12),
	.w2(32'h3a5edcee),
	.w3(32'hb97f280b),
	.w4(32'h39aea786),
	.w5(32'h3a95f35c),
	.w6(32'hbc2321b8),
	.w7(32'hbbdf2a22),
	.w8(32'hbc03d189),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc00ff92),
	.w1(32'hba99b79a),
	.w2(32'hbc28aee6),
	.w3(32'h39e23d15),
	.w4(32'h3adaf815),
	.w5(32'hbbaa4536),
	.w6(32'hba85d1d6),
	.w7(32'hba8002e1),
	.w8(32'hba18e075),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbef21d6),
	.w1(32'hbc0c2ed2),
	.w2(32'hbc26b5d0),
	.w3(32'hbc352a8b),
	.w4(32'hbbb3f5d5),
	.w5(32'hbbbbeb85),
	.w6(32'hbc1ad8d3),
	.w7(32'hbc081931),
	.w8(32'hbc34f9fc),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe6ab9b),
	.w1(32'hbc4da946),
	.w2(32'hbc9873b7),
	.w3(32'hbbe8278b),
	.w4(32'hbc13d18a),
	.w5(32'hbc347a43),
	.w6(32'hbbc72539),
	.w7(32'hbbd540f4),
	.w8(32'hbbcedab2),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6fd42c),
	.w1(32'hbb536373),
	.w2(32'hbbd9883a),
	.w3(32'hbb18e0c8),
	.w4(32'hba035e35),
	.w5(32'hbb0e05e0),
	.w6(32'hbbeed0b2),
	.w7(32'hbbf8bbc9),
	.w8(32'hbbedbb88),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd58515),
	.w1(32'hbba8b2b7),
	.w2(32'hbc1b51d5),
	.w3(32'hbb0fb262),
	.w4(32'hbb42775b),
	.w5(32'hbba10b9e),
	.w6(32'hbb07ec37),
	.w7(32'hbb6760d4),
	.w8(32'hbb111a05),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb393d8),
	.w1(32'hbbe75a0c),
	.w2(32'hbb8bb108),
	.w3(32'hbac00c0b),
	.w4(32'hbbc8160e),
	.w5(32'hbbe5319e),
	.w6(32'hbc1f1823),
	.w7(32'hbb94d9c7),
	.w8(32'hbc5d8f22),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc7ad57),
	.w1(32'hbb861833),
	.w2(32'hbabf1d4e),
	.w3(32'hbbb70cb8),
	.w4(32'hbbc6114d),
	.w5(32'hbbc8e5be),
	.w6(32'hba7be421),
	.w7(32'h3aa19fca),
	.w8(32'hbb03264f),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb915caaf),
	.w1(32'hbbd2787e),
	.w2(32'hbbfacce7),
	.w3(32'hbb8c4bcc),
	.w4(32'hbc2b640d),
	.w5(32'hbc64759e),
	.w6(32'hbbfd8b54),
	.w7(32'hbac8f639),
	.w8(32'hbc1229e5),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbde8841),
	.w1(32'hb91fa40d),
	.w2(32'hbaac0f6c),
	.w3(32'hbbe673d1),
	.w4(32'h3a8b847f),
	.w5(32'h3aa7aa3e),
	.w6(32'h3a3e361e),
	.w7(32'h3ae224cc),
	.w8(32'h3a342a65),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c002f9d),
	.w1(32'hbbb6ce96),
	.w2(32'hbc70872c),
	.w3(32'h3b5f7f6d),
	.w4(32'hbc18d90e),
	.w5(32'hbc59ae69),
	.w6(32'hbca5f0e2),
	.w7(32'hbcb31a91),
	.w8(32'hbcabefab),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc87e1d7),
	.w1(32'hbc101a3a),
	.w2(32'hbbbc3f7d),
	.w3(32'hbc313271),
	.w4(32'hbc036dbf),
	.w5(32'hbc816ddf),
	.w6(32'hbba75ef5),
	.w7(32'h3b977f62),
	.w8(32'h39a1b2cf),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4e8d2c),
	.w1(32'hbbaa8bb4),
	.w2(32'hbc00df00),
	.w3(32'hbbcda02c),
	.w4(32'hbba325de),
	.w5(32'hbbea914e),
	.w6(32'hbb6cd764),
	.w7(32'hbbca7b14),
	.w8(32'hbb033f41),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb598b5e),
	.w1(32'h3b8efcae),
	.w2(32'hbbe8f9ae),
	.w3(32'hbb4b5573),
	.w4(32'h3b63c3a4),
	.w5(32'hbbe6ed1b),
	.w6(32'h3c082bee),
	.w7(32'h39940a9a),
	.w8(32'h3b8cbbb5),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6f5d6d),
	.w1(32'hbbc75da1),
	.w2(32'hb9c28c60),
	.w3(32'hb908cd28),
	.w4(32'hbb654af2),
	.w5(32'h380bbfc8),
	.w6(32'hbbdb03cc),
	.w7(32'hbb5bc645),
	.w8(32'hbb924c16),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3cf212),
	.w1(32'hbb52b029),
	.w2(32'hbbbc6241),
	.w3(32'hba1bee8f),
	.w4(32'h39ad8eb7),
	.w5(32'hbb3bbf94),
	.w6(32'hbb9b4bdc),
	.w7(32'hbbd87a99),
	.w8(32'hbbdbcaf2),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaacfb0),
	.w1(32'hbb0f62e7),
	.w2(32'hbbe44c0a),
	.w3(32'h398880f0),
	.w4(32'h3b06bb54),
	.w5(32'hbb1f4e34),
	.w6(32'hbaa7cfd2),
	.w7(32'h3af2195b),
	.w8(32'hb8048786),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8af980),
	.w1(32'h3999321c),
	.w2(32'hb881e830),
	.w3(32'hb9af4cb4),
	.w4(32'hbb2902f9),
	.w5(32'hbb8c3faa),
	.w6(32'hba9ecd00),
	.w7(32'hbaf664e7),
	.w8(32'hbb4749e9),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdb00bc),
	.w1(32'hbc463822),
	.w2(32'hbc6d142a),
	.w3(32'hbbcad4ec),
	.w4(32'hbb00ee37),
	.w5(32'h3b95336f),
	.w6(32'hbc183c32),
	.w7(32'hbbc83331),
	.w8(32'hbbc6aab0),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbed4290),
	.w1(32'hba516f86),
	.w2(32'hbb87b9f9),
	.w3(32'h3988deff),
	.w4(32'h3a359d23),
	.w5(32'hbbf802e3),
	.w6(32'hbb02e1cd),
	.w7(32'hbb668367),
	.w8(32'hbb9a049d),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc177bde),
	.w1(32'hbbd50df0),
	.w2(32'hbc399a4f),
	.w3(32'hbbcda2af),
	.w4(32'hbb83cb6f),
	.w5(32'hbb7c1bac),
	.w6(32'hbb4c59ba),
	.w7(32'hbb94ebb7),
	.w8(32'hbb8fb762),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b018eb1),
	.w1(32'hb99ab7ed),
	.w2(32'hbc06e363),
	.w3(32'h3a394363),
	.w4(32'hbb098d49),
	.w5(32'hbc354ab1),
	.w6(32'hbb248ee7),
	.w7(32'hb9610ca7),
	.w8(32'hbbc9063c),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc01608b),
	.w1(32'hbbc4e993),
	.w2(32'hbbbb63d2),
	.w3(32'hbbf8fcdf),
	.w4(32'hbbc343bc),
	.w5(32'hbbe5730f),
	.w6(32'hbb05da4a),
	.w7(32'hbaef4fa3),
	.w8(32'hbbda7041),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad48a0a),
	.w1(32'h398bbef2),
	.w2(32'hba971563),
	.w3(32'h3b2ca589),
	.w4(32'h39bceb3a),
	.w5(32'h39621ca5),
	.w6(32'h3a26247e),
	.w7(32'hba0356c2),
	.w8(32'h3a963535),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aab0107),
	.w1(32'h3c16e77f),
	.w2(32'h3b87c5e6),
	.w3(32'h3b36ca52),
	.w4(32'h3c311358),
	.w5(32'h3bd8026f),
	.w6(32'h3c212b63),
	.w7(32'h3bd2f1fd),
	.w8(32'h3b51411e),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7b7622),
	.w1(32'h3c02744c),
	.w2(32'hbaa011b3),
	.w3(32'h3ba3de10),
	.w4(32'h3bd0509c),
	.w5(32'hbb24f9d0),
	.w6(32'h3b4addfb),
	.w7(32'hbab0222e),
	.w8(32'hbbdb0d60),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac84cb8),
	.w1(32'h3bf005be),
	.w2(32'hbb498a50),
	.w3(32'hbb54fd07),
	.w4(32'h3bcdadfa),
	.w5(32'hbba93128),
	.w6(32'h3b51d33e),
	.w7(32'hbb228596),
	.w8(32'hba71de7c),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb73dfc5),
	.w1(32'h397ef025),
	.w2(32'hbaa16c61),
	.w3(32'hbb951f95),
	.w4(32'hbac44406),
	.w5(32'hbb178e7a),
	.w6(32'h3808f752),
	.w7(32'hba864f02),
	.w8(32'hbad6791d),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba54c8cd),
	.w1(32'hba0f6e80),
	.w2(32'hbad1800f),
	.w3(32'hbabd2632),
	.w4(32'hb94c31d9),
	.w5(32'hba460817),
	.w6(32'hb99ab5a9),
	.w7(32'hba972705),
	.w8(32'h36a193df),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3543b0),
	.w1(32'h3b38a380),
	.w2(32'hbb415bf6),
	.w3(32'hb866236a),
	.w4(32'h3a4f5998),
	.w5(32'h3b0e8bab),
	.w6(32'h3ae98d66),
	.w7(32'h392a9bb2),
	.w8(32'h3add701b),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be03d1a),
	.w1(32'h3bb26fc4),
	.w2(32'hbbc7c243),
	.w3(32'h3c333d6d),
	.w4(32'h3c1f3aab),
	.w5(32'hbb195ef5),
	.w6(32'h3bebf674),
	.w7(32'h3a4bf49a),
	.w8(32'h3c551437),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8639f9),
	.w1(32'h3c1e32e2),
	.w2(32'h3c5c9db5),
	.w3(32'h3c336484),
	.w4(32'h3bfb3abb),
	.w5(32'h3c06b823),
	.w6(32'h3aa904ab),
	.w7(32'h3bdf960f),
	.w8(32'h3b619b79),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c188485),
	.w1(32'hba07657e),
	.w2(32'hbb23931e),
	.w3(32'h3c00438a),
	.w4(32'hbaf604e3),
	.w5(32'hbb3c55b6),
	.w6(32'hbb103bc1),
	.w7(32'hbb5ea556),
	.w8(32'hbb36e4c0),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafb82ef),
	.w1(32'h3b34b1f1),
	.w2(32'h3bc78e0c),
	.w3(32'hba95143f),
	.w4(32'h3ae5668b),
	.w5(32'h3b474e50),
	.w6(32'h3ac7c459),
	.w7(32'h3b06808f),
	.w8(32'hbae15364),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad13405),
	.w1(32'hbc7069dd),
	.w2(32'hbc6f96e1),
	.w3(32'h3ade0869),
	.w4(32'hbc2f4076),
	.w5(32'hbc18ab78),
	.w6(32'hbc390856),
	.w7(32'hbc3a7b6c),
	.w8(32'hbbde985e),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0c53f7),
	.w1(32'hbb54afac),
	.w2(32'hbbacf422),
	.w3(32'hbbd0ad86),
	.w4(32'hb98211f2),
	.w5(32'hba46d2fe),
	.w6(32'hbae26a4d),
	.w7(32'hbb53b0f3),
	.w8(32'h39bc82a4),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b08bd60),
	.w1(32'hbb9602be),
	.w2(32'hbc033d71),
	.w3(32'h3b480a0f),
	.w4(32'hba9ec9fe),
	.w5(32'hbb68bff0),
	.w6(32'hbbbdba3d),
	.w7(32'hbbd3012d),
	.w8(32'hbbae3eb8),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb3b847),
	.w1(32'hbada34f3),
	.w2(32'hbc2233e1),
	.w3(32'hba77c586),
	.w4(32'hbb225e06),
	.w5(32'hbc52ee54),
	.w6(32'hbb15fa53),
	.w7(32'hbc093b5b),
	.w8(32'hbc0a3a17),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc6de6e),
	.w1(32'h3aab9aae),
	.w2(32'h3b1919fe),
	.w3(32'hbc01dda4),
	.w4(32'hbb383b20),
	.w5(32'hbb1f79b0),
	.w6(32'h37194e71),
	.w7(32'hba6c3f6a),
	.w8(32'hbb077010),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a887d22),
	.w1(32'hb8840975),
	.w2(32'hbbb8a1a1),
	.w3(32'h3aaea89a),
	.w4(32'h3a905002),
	.w5(32'hbb39eb25),
	.w6(32'hbb425d00),
	.w7(32'hbb3951f2),
	.w8(32'hbb6c0363),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9905476),
	.w1(32'hbbe881b6),
	.w2(32'hbb5ac0aa),
	.w3(32'hbabdc793),
	.w4(32'hbc4f306a),
	.w5(32'hbc1914e0),
	.w6(32'hbc61afe1),
	.w7(32'hbc093db0),
	.w8(32'hbca52225),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbdacdd),
	.w1(32'hbbcd8253),
	.w2(32'hbc8e906b),
	.w3(32'hbcac4579),
	.w4(32'h3b4dcb47),
	.w5(32'hbb049342),
	.w6(32'hbbb6cc74),
	.w7(32'h38c50fe9),
	.w8(32'hbb0eb50a),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3fe362),
	.w1(32'hbb86da82),
	.w2(32'hbc29cbe0),
	.w3(32'hbb581e3f),
	.w4(32'h3b904563),
	.w5(32'h3b9a0a18),
	.w6(32'hba22b84e),
	.w7(32'hbaab05da),
	.w8(32'h3b57ae65),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h382e6c17),
	.w1(32'hbc0083a3),
	.w2(32'hbc5840c2),
	.w3(32'h3bc346e9),
	.w4(32'hbc239e12),
	.w5(32'hbc64c01f),
	.w6(32'hbbbc18fa),
	.w7(32'h3a9de8af),
	.w8(32'hbb890469),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb030611),
	.w1(32'h3c0784c9),
	.w2(32'h3adfd937),
	.w3(32'hbb2c0c00),
	.w4(32'h3ba1a86b),
	.w5(32'hba883b5d),
	.w6(32'h3c06ad91),
	.w7(32'h3ac5f20a),
	.w8(32'h3b04de94),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb83cb32),
	.w1(32'hbb916578),
	.w2(32'hbc1342dd),
	.w3(32'hbb6c2d11),
	.w4(32'hbb4148e8),
	.w5(32'hbb972cb8),
	.w6(32'hbb8a9bfe),
	.w7(32'hbb69ac07),
	.w8(32'hbb1f2269),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba159716),
	.w1(32'hbc21577f),
	.w2(32'hbc3bf1d6),
	.w3(32'h392071f3),
	.w4(32'hbbbd65d5),
	.w5(32'hbbbd4fc9),
	.w6(32'hbc0c9805),
	.w7(32'hbc164c45),
	.w8(32'hbbe7ae2e),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd934a3),
	.w1(32'hbc567d61),
	.w2(32'hbc73fd00),
	.w3(32'hbb9e9c7d),
	.w4(32'hbc02d759),
	.w5(32'hbc19048b),
	.w6(32'hbc45c601),
	.w7(32'hbc34c3c7),
	.w8(32'hbbcad56d),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b3b14),
	.w1(32'h39d18efb),
	.w2(32'hbc3d7ac2),
	.w3(32'hbb0956a2),
	.w4(32'hbbcd9f9f),
	.w5(32'hbc83e4fb),
	.w6(32'hb721e1e3),
	.w7(32'hbbb86769),
	.w8(32'hbc597a0b),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbcc989),
	.w1(32'hbc4c6f67),
	.w2(32'hbc94799e),
	.w3(32'hbc9aac21),
	.w4(32'hbc797015),
	.w5(32'hbc863b02),
	.w6(32'hbc93d18a),
	.w7(32'hbc8c9bf5),
	.w8(32'hbc82b201),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6008da),
	.w1(32'h39bdfc36),
	.w2(32'hbbaa7860),
	.w3(32'hbc6b318b),
	.w4(32'h39e7eb5b),
	.w5(32'hbb887ae9),
	.w6(32'hb9aab4c7),
	.w7(32'hbb998136),
	.w8(32'hbb94e8e4),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d6c3e),
	.w1(32'hba9c3c63),
	.w2(32'hbad23a70),
	.w3(32'hbba6b8fb),
	.w4(32'hbba0f79a),
	.w5(32'hbbbec3de),
	.w6(32'hbb592ca9),
	.w7(32'hbba77d0c),
	.w8(32'hbb718a26),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1d210f),
	.w1(32'h3be1beb8),
	.w2(32'h3ab22263),
	.w3(32'hbb4faa8d),
	.w4(32'h3b2f2c07),
	.w5(32'hbb6f10e9),
	.w6(32'hba88b7b3),
	.w7(32'hbafe620f),
	.w8(32'hbbd9fc2a),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc37a9ce),
	.w1(32'hbc19674f),
	.w2(32'hbc5886e0),
	.w3(32'hbc40e8b4),
	.w4(32'hbbf6ddf0),
	.w5(32'hbc674c3d),
	.w6(32'hbbc0acfc),
	.w7(32'hbc3637c6),
	.w8(32'hbc3b75c4),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc55507c),
	.w1(32'hbc73e751),
	.w2(32'hbc5b88dd),
	.w3(32'hbc357638),
	.w4(32'hbc0165bc),
	.w5(32'hbc0906cc),
	.w6(32'hbba3ce20),
	.w7(32'hbc140bf4),
	.w8(32'hbb99d1fe),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b37ec33),
	.w1(32'hbc04a1f2),
	.w2(32'hbc20d332),
	.w3(32'hbb4e7602),
	.w4(32'hbb26ea7b),
	.w5(32'hbb6f3106),
	.w6(32'hbbef3739),
	.w7(32'hbc054677),
	.w8(32'hbb88f1ae),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc82240d),
	.w1(32'hbbcf3927),
	.w2(32'hbc81434a),
	.w3(32'hbb20f96f),
	.w4(32'h3ba4dc0e),
	.w5(32'hb8ac5228),
	.w6(32'hbafbde8b),
	.w7(32'h3bb37e38),
	.w8(32'h3b031ebd),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3983aa36),
	.w1(32'hbc14d4a2),
	.w2(32'hbc91d31d),
	.w3(32'hb9fad6f7),
	.w4(32'hbb53f62e),
	.w5(32'hbc219bf0),
	.w6(32'hbc2cb7a4),
	.w7(32'hbc0d9915),
	.w8(32'hbc630e09),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdc58b1),
	.w1(32'hbbdf5d76),
	.w2(32'hbbf867d0),
	.w3(32'hbb63bf75),
	.w4(32'hbbb9f64e),
	.w5(32'hbb856d5c),
	.w6(32'hbb55a0ce),
	.w7(32'hbba6ac39),
	.w8(32'hbb72240e),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb99658d),
	.w1(32'hbb749c9f),
	.w2(32'hbb70bd2b),
	.w3(32'hbb05f052),
	.w4(32'hbb76d8d8),
	.w5(32'hbb1c0b9d),
	.w6(32'hbc1fa330),
	.w7(32'hbba9cadf),
	.w8(32'h3b209055),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb08b14c),
	.w1(32'hbb4152d2),
	.w2(32'h3a77154f),
	.w3(32'hbac1b91c),
	.w4(32'hbbd5086d),
	.w5(32'hbb844da9),
	.w6(32'hbbdda63b),
	.w7(32'hbb92fbee),
	.w8(32'hbc3f3bc0),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc16a38b),
	.w1(32'h3a0c9ccf),
	.w2(32'h3b9d3d2e),
	.w3(32'hbc2235bf),
	.w4(32'h3b256181),
	.w5(32'h3b93756a),
	.w6(32'h3aa5e9d2),
	.w7(32'h3b9213fb),
	.w8(32'h3b9584a5),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bae0029),
	.w1(32'hbb26a028),
	.w2(32'hbc0c46d6),
	.w3(32'h3be3c9ad),
	.w4(32'hbaa5904a),
	.w5(32'hbb973b76),
	.w6(32'h3b49f71f),
	.w7(32'hbbc9dea2),
	.w8(32'hba3f67aa),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0b46e9),
	.w1(32'h3bc35bf3),
	.w2(32'hb9262dff),
	.w3(32'h3bb359db),
	.w4(32'h3c02d9a8),
	.w5(32'h3ac2b8a5),
	.w6(32'h3be2c651),
	.w7(32'h3bb7338f),
	.w8(32'hba920c52),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0aa765),
	.w1(32'h3b1aadeb),
	.w2(32'hbb6a288d),
	.w3(32'h3a8c67c7),
	.w4(32'h3ba1bdc4),
	.w5(32'hbbefca3b),
	.w6(32'h39bd6345),
	.w7(32'hbb452716),
	.w8(32'hbb759b18),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7ef34f),
	.w1(32'hbb45ca49),
	.w2(32'hbbc83899),
	.w3(32'hbb8acf2c),
	.w4(32'hbb788907),
	.w5(32'hbbcac266),
	.w6(32'hbb627d6c),
	.w7(32'hbbcf184f),
	.w8(32'hbb8ab3d6),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe3698e),
	.w1(32'hbba91826),
	.w2(32'hbc00e981),
	.w3(32'hbabc25c5),
	.w4(32'h3bc23d3f),
	.w5(32'h3b964ac8),
	.w6(32'hbb15133d),
	.w7(32'h3b1c1bf4),
	.w8(32'h3a9d5eb4),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbeb83d),
	.w1(32'hbbb3b8de),
	.w2(32'hbb4e7b5a),
	.w3(32'h3be94d6d),
	.w4(32'hbb9546cf),
	.w5(32'hbb283cb7),
	.w6(32'hbac1d36c),
	.w7(32'hbb1e2306),
	.w8(32'hbb09966c),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbace2262),
	.w1(32'hbae196ba),
	.w2(32'hbb7fe20f),
	.w3(32'h39cf014d),
	.w4(32'hba4f85a4),
	.w5(32'hba9de967),
	.w6(32'hba8b57be),
	.w7(32'hbb35dab1),
	.w8(32'hbb03f14c),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0602ae),
	.w1(32'hbbbb8e74),
	.w2(32'hbba97491),
	.w3(32'hbb95b38f),
	.w4(32'hbae9b0bf),
	.w5(32'hb7a8f4e4),
	.w6(32'hbb8d4695),
	.w7(32'hbb79da67),
	.w8(32'hb8a0cd2a),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398189fe),
	.w1(32'hba5dc13a),
	.w2(32'hbb2f1573),
	.w3(32'h3af08081),
	.w4(32'hbae7ccfe),
	.w5(32'hbb345e92),
	.w6(32'hba811bcc),
	.w7(32'hbb38f63a),
	.w8(32'hbabfc4fb),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3d1d2c),
	.w1(32'hbb5ed2c4),
	.w2(32'hbba4694d),
	.w3(32'h3a15c780),
	.w4(32'hbac84f52),
	.w5(32'hbb590552),
	.w6(32'hbb4835ff),
	.w7(32'hbb716576),
	.w8(32'hba5b1ed3),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbba7a49),
	.w1(32'h3b926090),
	.w2(32'hbb2350a2),
	.w3(32'hbba8614c),
	.w4(32'hbc39126b),
	.w5(32'hbca10f07),
	.w6(32'h3a01b4e4),
	.w7(32'h3aadaa7e),
	.w8(32'hbc962794),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3acf35),
	.w1(32'hbb94da07),
	.w2(32'hbbc3ce59),
	.w3(32'hbc16390b),
	.w4(32'hbb137a77),
	.w5(32'hbb24a4bb),
	.w6(32'hbc195043),
	.w7(32'hbc00ac0c),
	.w8(32'hbc30d83a),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb804c10),
	.w1(32'hbb9c3fcb),
	.w2(32'hbbb31bb2),
	.w3(32'hbb96e676),
	.w4(32'hbb8fe600),
	.w5(32'hbb8c30c8),
	.w6(32'hbbe1e111),
	.w7(32'hbbed4c92),
	.w8(32'hbba25597),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc97b64),
	.w1(32'h3c0f673f),
	.w2(32'h3a316196),
	.w3(32'hbb2c9ca7),
	.w4(32'h3a4410fc),
	.w5(32'hbbf7cb7a),
	.w6(32'h3bb18039),
	.w7(32'hb99c93c1),
	.w8(32'hbba29e1e),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1c4977),
	.w1(32'h3b410b88),
	.w2(32'h3afe3911),
	.w3(32'hbb092c14),
	.w4(32'h3b37b660),
	.w5(32'h3b3f24b8),
	.w6(32'hb8c501f9),
	.w7(32'h3b75c3ca),
	.w8(32'h39d28366),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7bacba),
	.w1(32'h3c0c4030),
	.w2(32'h3a3483c2),
	.w3(32'h3a336bed),
	.w4(32'h3c2f90e8),
	.w5(32'h39d449bd),
	.w6(32'h3bbc353c),
	.w7(32'h3be78cab),
	.w8(32'h3a571e37),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a02de5c),
	.w1(32'h3b06d576),
	.w2(32'h3b7d6cd3),
	.w3(32'hbb15c2f9),
	.w4(32'h3b0c1ae5),
	.w5(32'h3b7202c8),
	.w6(32'h3afd096f),
	.w7(32'h3b61a4c4),
	.w8(32'h3b44103d),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4ce583),
	.w1(32'hbaa8c433),
	.w2(32'hbb84cd23),
	.w3(32'h3b74f88e),
	.w4(32'hbb91f275),
	.w5(32'hbc021e77),
	.w6(32'hbb7d7c70),
	.w7(32'hbbc8e61c),
	.w8(32'hbbedade2),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc45a2e5),
	.w1(32'hbc3f0d7f),
	.w2(32'hbc660cca),
	.w3(32'hbb998fe3),
	.w4(32'hbb6102c1),
	.w5(32'hbbce2457),
	.w6(32'hbba5521d),
	.w7(32'hbc16342a),
	.w8(32'hbc27319f),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc234a08),
	.w1(32'hbb634645),
	.w2(32'hbbf4bc88),
	.w3(32'hbad9d96e),
	.w4(32'h3a8061c8),
	.w5(32'hbc06e794),
	.w6(32'hbb1b8d23),
	.w7(32'hbbaeffe8),
	.w8(32'hbb615987),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb627e96),
	.w1(32'hb9dd866d),
	.w2(32'hbbc246d4),
	.w3(32'h39b8653a),
	.w4(32'h3b4f6b78),
	.w5(32'hbafca35d),
	.w6(32'hb99be9ab),
	.w7(32'h3a1508f1),
	.w8(32'hbbb2a4d1),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a9036),
	.w1(32'h3bd525ab),
	.w2(32'h3b87605c),
	.w3(32'hbbd25874),
	.w4(32'hbaa671a6),
	.w5(32'hba1c4a7e),
	.w6(32'h3b3974ad),
	.w7(32'h3a665da3),
	.w8(32'hba3c51ee),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5de466),
	.w1(32'h3a523a65),
	.w2(32'h3a0f1290),
	.w3(32'h3b1e43be),
	.w4(32'hb9cbdd43),
	.w5(32'hba348207),
	.w6(32'h39c273f2),
	.w7(32'hb97ca897),
	.w8(32'h39c2a58c),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0ca21f),
	.w1(32'hbc4688e4),
	.w2(32'hbc3c53b9),
	.w3(32'hbb0291a1),
	.w4(32'hbc465aa3),
	.w5(32'hbc4cb2e1),
	.w6(32'hbc4d54b7),
	.w7(32'hbc5d0aba),
	.w8(32'hbc1de9c1),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc30ae5d),
	.w1(32'hbb726644),
	.w2(32'hbb2e7796),
	.w3(32'hbc22e016),
	.w4(32'hbbfc4d6c),
	.w5(32'hbbe4a011),
	.w6(32'h3b84b008),
	.w7(32'hbb09735e),
	.w8(32'hbb976b49),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdf2c03),
	.w1(32'hb9e5be9f),
	.w2(32'hbbb37056),
	.w3(32'hba808bac),
	.w4(32'h3b3e755a),
	.w5(32'hbae1582e),
	.w6(32'hbac5b424),
	.w7(32'h3b3b6582),
	.w8(32'h39dcb6a3),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb97fa55),
	.w1(32'hbc511060),
	.w2(32'hbc17de55),
	.w3(32'hbaf53a7e),
	.w4(32'hbc5ef0d4),
	.w5(32'hbc2c6949),
	.w6(32'hbc30b44b),
	.w7(32'hbc1b448d),
	.w8(32'hbc6d999b),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc11af82),
	.w1(32'h3c0f644c),
	.w2(32'h3c243589),
	.w3(32'hbc4604d8),
	.w4(32'h3b814584),
	.w5(32'h3b0650c7),
	.w6(32'hb98af687),
	.w7(32'h3b0ed2f3),
	.w8(32'hbb1a7603),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4b3e8f),
	.w1(32'h3bebe521),
	.w2(32'hb9f6ef1e),
	.w3(32'hbb1a171a),
	.w4(32'h3bbccf45),
	.w5(32'hbb8a02cc),
	.w6(32'h3a403ae5),
	.w7(32'h37fecd13),
	.w8(32'hbc07792c),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad5856f),
	.w1(32'hbb9fb906),
	.w2(32'hbb6d0d0a),
	.w3(32'hbb53b7e0),
	.w4(32'hbb1432d0),
	.w5(32'hbacf0dc7),
	.w6(32'hbb822d79),
	.w7(32'hbb97d51a),
	.w8(32'hbb025075),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4a99e9),
	.w1(32'hbc0d8911),
	.w2(32'hbc1e0854),
	.w3(32'hbada7626),
	.w4(32'hbc127e15),
	.w5(32'hbbd86d51),
	.w6(32'hbbba652a),
	.w7(32'hbbd36516),
	.w8(32'hbbaefed2),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc33f18),
	.w1(32'hbbb9cfe6),
	.w2(32'hb99a69ee),
	.w3(32'hbb7d29ef),
	.w4(32'hbbcbb1ac),
	.w5(32'hbb9a1276),
	.w6(32'hbbf2cbf4),
	.w7(32'hbbbe0774),
	.w8(32'hbbc2bef0),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc5c3d1),
	.w1(32'hbb319b9f),
	.w2(32'h3a579ffd),
	.w3(32'hbbada0dd),
	.w4(32'hba85c1b2),
	.w5(32'h3b2754cc),
	.w6(32'hbadc205f),
	.w7(32'h3a653b3a),
	.w8(32'h3b956168),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba0d630),
	.w1(32'hbc055c49),
	.w2(32'hbc0281f2),
	.w3(32'h3b8bd47e),
	.w4(32'hbbbd6f7a),
	.w5(32'hbbb7ec3d),
	.w6(32'hbb40f67f),
	.w7(32'hbbb64dc5),
	.w8(32'hbb2d738f),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe793d1),
	.w1(32'h3b17c4d6),
	.w2(32'h3b0d398a),
	.w3(32'hb9feabcf),
	.w4(32'h3a81bd40),
	.w5(32'hbb54c34b),
	.w6(32'hb9b194e7),
	.w7(32'hbb8dbbf1),
	.w8(32'hbb901c45),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3435f5),
	.w1(32'hbbfea622),
	.w2(32'hbb84a2b5),
	.w3(32'h3a91daa2),
	.w4(32'hba813504),
	.w5(32'hbb24f0bf),
	.w6(32'hbbc1249e),
	.w7(32'hbba648e4),
	.w8(32'hbb8165f9),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c083bca),
	.w1(32'hbb0223cd),
	.w2(32'hbc5e863b),
	.w3(32'hba6c699a),
	.w4(32'hba183fb0),
	.w5(32'hbbc5b0a7),
	.w6(32'h3aed1244),
	.w7(32'hbbde5701),
	.w8(32'hba8e4930),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc81411f),
	.w1(32'hbc520cc2),
	.w2(32'hbc4d37aa),
	.w3(32'hbb73f162),
	.w4(32'hbbfe2e25),
	.w5(32'hbb91bacd),
	.w6(32'hbc2c799c),
	.w7(32'hbc2ec3f6),
	.w8(32'hbc5491fe),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe56249),
	.w1(32'hbb926864),
	.w2(32'hbbc5de7e),
	.w3(32'hbbafbc02),
	.w4(32'hba8fdcbc),
	.w5(32'hba88ba01),
	.w6(32'hbb725ee1),
	.w7(32'hbb647bcf),
	.w8(32'hbb31226a),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae9d6ee),
	.w1(32'hbb204186),
	.w2(32'hbac0fee0),
	.w3(32'hba2dce83),
	.w4(32'hbb06a3be),
	.w5(32'hb9ad691b),
	.w6(32'hbb97f1c3),
	.w7(32'hbb87059a),
	.w8(32'hbb8fffc8),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb764b74),
	.w1(32'hba7a951a),
	.w2(32'hbb688e1b),
	.w3(32'hbb42d2ba),
	.w4(32'hba633b98),
	.w5(32'hba5e9f49),
	.w6(32'hb9dd1942),
	.w7(32'hb9e72196),
	.w8(32'h3a3f891b),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c46af7),
	.w1(32'hbb790d9a),
	.w2(32'hbb14310a),
	.w3(32'h3a9d65a8),
	.w4(32'hba88f542),
	.w5(32'hb99cd952),
	.w6(32'hbb77bd63),
	.w7(32'hbb70a7dc),
	.w8(32'hbac011a5),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb02be2a),
	.w1(32'h396620ae),
	.w2(32'hba615fbe),
	.w3(32'hba38dd10),
	.w4(32'hbb3077cd),
	.w5(32'hbb97534d),
	.w6(32'hbaa135a2),
	.w7(32'hbb2571de),
	.w8(32'hbaa7e20c),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae51c4f),
	.w1(32'hbb841b04),
	.w2(32'hbb579781),
	.w3(32'hbb4a39bd),
	.w4(32'hbb3279a1),
	.w5(32'hba548ff4),
	.w6(32'hbbc4df22),
	.w7(32'hbbb86cc0),
	.w8(32'hbbacf13d),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb265898),
	.w1(32'hbbc55712),
	.w2(32'hbc0ef01c),
	.w3(32'hbb3cb9c7),
	.w4(32'hbb2bc66f),
	.w5(32'hbb309c2e),
	.w6(32'hbc11bad2),
	.w7(32'hbbee2bf2),
	.w8(32'hbb09a83b),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba89cb3),
	.w1(32'hbaff24b2),
	.w2(32'hbbdd1910),
	.w3(32'h3b0a120e),
	.w4(32'hba46421a),
	.w5(32'hbb926a7c),
	.w6(32'hbae5834c),
	.w7(32'hbb6f2031),
	.w8(32'hbaeb765c),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba26fcf),
	.w1(32'h3b4d459e),
	.w2(32'hbc5e9559),
	.w3(32'hbbc48563),
	.w4(32'hbb7da590),
	.w5(32'hbc4827e7),
	.w6(32'hbafec1c6),
	.w7(32'hba9c7929),
	.w8(32'hbc1810a6),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8b726d),
	.w1(32'hbbc2eafd),
	.w2(32'hbc602b54),
	.w3(32'hbc19073d),
	.w4(32'hbb184ddc),
	.w5(32'hbc00e91e),
	.w6(32'hbb51a3cf),
	.w7(32'hbb8efc27),
	.w8(32'hbb535f5f),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbffa2b9),
	.w1(32'hbba5a364),
	.w2(32'hbc01c548),
	.w3(32'hbb8588a6),
	.w4(32'hbb0db7b5),
	.w5(32'hbb8698b5),
	.w6(32'hbb5dcc2f),
	.w7(32'h3a441ce7),
	.w8(32'h3b052c39),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa46c54),
	.w1(32'h3bef266a),
	.w2(32'h3b761a6f),
	.w3(32'h3b3e28e1),
	.w4(32'h3bd09100),
	.w5(32'h3bb69f70),
	.w6(32'h3bde99fb),
	.w7(32'h3b8c49ce),
	.w8(32'h3bfff4e7),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb5b6d0),
	.w1(32'hbbbed1e3),
	.w2(32'hbb8639e9),
	.w3(32'h3c0a8ee2),
	.w4(32'hbb7f2b92),
	.w5(32'hba533c7a),
	.w6(32'hbc0c0b9a),
	.w7(32'hbbfcde6e),
	.w8(32'hbbf63b0a),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5c7686),
	.w1(32'hbae5ae02),
	.w2(32'hba2e11c6),
	.w3(32'hbb836e90),
	.w4(32'hbb213499),
	.w5(32'hba8ea6d9),
	.w6(32'hbab018a8),
	.w7(32'hbaa24ce0),
	.w8(32'hbad39f91),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a253e9e),
	.w1(32'h3a29e8f7),
	.w2(32'h3b100a0f),
	.w3(32'hba75e8e2),
	.w4(32'hb9f023b7),
	.w5(32'h3a54b138),
	.w6(32'hba22511e),
	.w7(32'hb9978734),
	.w8(32'hbae80d2d),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb8d0d6),
	.w1(32'hbc15d1e3),
	.w2(32'hbc3963e2),
	.w3(32'hbb874ead),
	.w4(32'hbafaced1),
	.w5(32'h3ae38c6c),
	.w6(32'hbc157e13),
	.w7(32'hbb89c8cc),
	.w8(32'hbb73c866),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9953ff),
	.w1(32'hbba88656),
	.w2(32'hbbf5111e),
	.w3(32'hbb22bfaf),
	.w4(32'hbaa1347c),
	.w5(32'hbb4dc0c5),
	.w6(32'hbb499c06),
	.w7(32'hbb919232),
	.w8(32'h3b4d3c02),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc2abf5),
	.w1(32'hbb1fc771),
	.w2(32'hbbda4fb6),
	.w3(32'h3b5333e6),
	.w4(32'hbaccfc68),
	.w5(32'hbb5da375),
	.w6(32'hbb6879e0),
	.w7(32'hbbda7586),
	.w8(32'hbbb4b6c0),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0525af),
	.w1(32'hbbb80f78),
	.w2(32'hbbfa6eca),
	.w3(32'hbbdff037),
	.w4(32'hbb83e5b4),
	.w5(32'hbbc2d8d0),
	.w6(32'hbb9347a9),
	.w7(32'hbbc04781),
	.w8(32'hbb353f24),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba5368f),
	.w1(32'hbb9f7c76),
	.w2(32'hbbe237a8),
	.w3(32'hbb81cda5),
	.w4(32'hbae7d370),
	.w5(32'hbae64320),
	.w6(32'hbb5ac26a),
	.w7(32'hbba72810),
	.w8(32'hbacc5d11),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb12d827),
	.w1(32'hbc4caffa),
	.w2(32'hbc5d487e),
	.w3(32'h3a9e590d),
	.w4(32'hbb0bedb0),
	.w5(32'hba3fad99),
	.w6(32'hbbe3856c),
	.w7(32'hbb1206fe),
	.w8(32'hba82c9ed),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc069eaf),
	.w1(32'hbb336e1b),
	.w2(32'hbb95cbf2),
	.w3(32'hbb93a2c9),
	.w4(32'hbbd92351),
	.w5(32'hbc0e38d7),
	.w6(32'hbb7c5069),
	.w7(32'hbbca5aea),
	.w8(32'hbba35f69),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2dadc4),
	.w1(32'h3a8e1493),
	.w2(32'hbbfd541a),
	.w3(32'hbc81d878),
	.w4(32'h3b635344),
	.w5(32'h3a9d24f4),
	.w6(32'hbb275bad),
	.w7(32'h3b782332),
	.w8(32'hbb4e0dfd),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaca5b13),
	.w1(32'hb90785b9),
	.w2(32'hb937b8e5),
	.w3(32'hbb1db686),
	.w4(32'hb8960abf),
	.w5(32'hb93014fe),
	.w6(32'h38649b9a),
	.w7(32'hb8c56df1),
	.w8(32'hb8a8f5eb),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a5a216),
	.w1(32'h39b62352),
	.w2(32'h392e42de),
	.w3(32'h3ab44823),
	.w4(32'h3b227fdc),
	.w5(32'hbab93d37),
	.w6(32'hbb00ea8d),
	.w7(32'hbaaf6504),
	.w8(32'hbb86d584),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule