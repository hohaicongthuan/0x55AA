module layer_10_featuremap_448(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba359742),
	.w1(32'h3b00f444),
	.w2(32'h386ec9d5),
	.w3(32'hbc1af75b),
	.w4(32'h3b81f4c8),
	.w5(32'hba03e5b7),
	.w6(32'hbacaf1a7),
	.w7(32'h3bfdd27e),
	.w8(32'h3c05d374),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc83dcb),
	.w1(32'h3ba488cd),
	.w2(32'h3ad6103b),
	.w3(32'hbc87a3db),
	.w4(32'h3c2db791),
	.w5(32'h3bc31ebf),
	.w6(32'hbba6ad65),
	.w7(32'h3c516579),
	.w8(32'h3a9e0ff7),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a7ba9a),
	.w1(32'hbb578340),
	.w2(32'hbc4a60d4),
	.w3(32'h3bac8e93),
	.w4(32'h3ca0aa84),
	.w5(32'hbc5c1d1d),
	.w6(32'h3bc21000),
	.w7(32'h3c3dcef6),
	.w8(32'h3d256937),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8f9073),
	.w1(32'hbc6f05e4),
	.w2(32'hbbc89eea),
	.w3(32'h3bd89d5c),
	.w4(32'hbc83c417),
	.w5(32'hbc4e2545),
	.w6(32'h3b472025),
	.w7(32'hbc9205f6),
	.w8(32'hbc21c75e),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc62386e),
	.w1(32'hbbe7f53d),
	.w2(32'hbbd00abc),
	.w3(32'hbc4ecf07),
	.w4(32'hbc630177),
	.w5(32'hbbe44875),
	.w6(32'hbbda7487),
	.w7(32'hbbc5aa9a),
	.w8(32'hbc817e52),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc0fb98),
	.w1(32'hbaeec265),
	.w2(32'h3c4013a6),
	.w3(32'h3b72afbc),
	.w4(32'hbc2f8bf4),
	.w5(32'h3b95cbde),
	.w6(32'hbc10c3ea),
	.w7(32'hbb6052b3),
	.w8(32'h3bc77384),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b46062c),
	.w1(32'hbae2deb7),
	.w2(32'hbc139479),
	.w3(32'h3bb1c5da),
	.w4(32'h3b078687),
	.w5(32'h3b36107f),
	.w6(32'h3be72973),
	.w7(32'hbb73a956),
	.w8(32'h3c33dddf),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c05788e),
	.w1(32'hbc2f1b10),
	.w2(32'hbd186981),
	.w3(32'h3c243148),
	.w4(32'h3c6b5d0f),
	.w5(32'h3c2f1c9e),
	.w6(32'hbc3ac625),
	.w7(32'h3af9a87a),
	.w8(32'h3d096387),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc87fabf),
	.w1(32'hbb272e2c),
	.w2(32'h3b7d2d05),
	.w3(32'hbc88d465),
	.w4(32'hbcb7333d),
	.w5(32'h3c5c1f15),
	.w6(32'hbc986af2),
	.w7(32'h3becc8d1),
	.w8(32'h3ce4467c),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd17925),
	.w1(32'h3b0d6ef9),
	.w2(32'h3bf8e5ad),
	.w3(32'h3d5efde2),
	.w4(32'hbb6cd3ed),
	.w5(32'hbc5434f5),
	.w6(32'h3a89fb1a),
	.w7(32'hbb18c68a),
	.w8(32'hbc20c536),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f896d5),
	.w1(32'hbb2ef7fc),
	.w2(32'hbaced848),
	.w3(32'hbbb01c0e),
	.w4(32'h399ae446),
	.w5(32'hbc35bbe1),
	.w6(32'h3bac179b),
	.w7(32'h3c37073f),
	.w8(32'h3b2462bf),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c16bde7),
	.w1(32'hbbd8378a),
	.w2(32'h3b27ee7f),
	.w3(32'h3c536c0f),
	.w4(32'hbcb2f84d),
	.w5(32'h3ba7d153),
	.w6(32'h3c1f7d1a),
	.w7(32'hbc1cc560),
	.w8(32'h3b254763),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c83040a),
	.w1(32'hbc51959e),
	.w2(32'h3b896b75),
	.w3(32'h3cbeab96),
	.w4(32'hbbbec19d),
	.w5(32'h3cb048ae),
	.w6(32'h3be8c73c),
	.w7(32'hbbb271b9),
	.w8(32'hbb4515d2),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd084a4),
	.w1(32'hbcd768f6),
	.w2(32'h3c6aac5e),
	.w3(32'hbc32f1a6),
	.w4(32'hbc9264c9),
	.w5(32'h3c5fcaef),
	.w6(32'hbc29ce5e),
	.w7(32'hbc0634cb),
	.w8(32'hbca55ac3),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcdec02a),
	.w1(32'hbb99d66e),
	.w2(32'hbbf19b89),
	.w3(32'hbc039952),
	.w4(32'hbb474228),
	.w5(32'hbc0d7eb8),
	.w6(32'hbbfb4667),
	.w7(32'hba7ce278),
	.w8(32'hbc69873f),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdac20d),
	.w1(32'h3b723329),
	.w2(32'hbbce9a65),
	.w3(32'hbc2ee45a),
	.w4(32'h3c07e5c6),
	.w5(32'hbb807dda),
	.w6(32'hbc3db390),
	.w7(32'h3b55fa37),
	.w8(32'hba80ae5b),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac4c0a3),
	.w1(32'h3bb748e4),
	.w2(32'h3b8a5ff4),
	.w3(32'hbbf98a35),
	.w4(32'h3a9da83c),
	.w5(32'h3a2086be),
	.w6(32'hbb533aad),
	.w7(32'hbb99a160),
	.w8(32'hbbf52f36),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab280b9),
	.w1(32'h3c29a704),
	.w2(32'h3a259eb1),
	.w3(32'hbb63040a),
	.w4(32'h3c53db25),
	.w5(32'hbc8c1175),
	.w6(32'hbc129f48),
	.w7(32'h3b380fed),
	.w8(32'hbc2bab67),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb563933),
	.w1(32'hb8e7eb7b),
	.w2(32'h3aebef58),
	.w3(32'hbd13c4df),
	.w4(32'hbc8e9bdb),
	.w5(32'h3ba81fd6),
	.w6(32'hbcda3503),
	.w7(32'hbb9735b9),
	.w8(32'h3bddf4c7),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b116acd),
	.w1(32'h3b5edbe0),
	.w2(32'h3ba4b1fe),
	.w3(32'h3d074008),
	.w4(32'h3acfb4c8),
	.w5(32'hbc6876c0),
	.w6(32'h3b950444),
	.w7(32'h3c24c904),
	.w8(32'hbb256192),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc00b0f),
	.w1(32'h3a3e81ed),
	.w2(32'h3a8819b2),
	.w3(32'h39c3a8bc),
	.w4(32'hbbe5aefb),
	.w5(32'h3b291820),
	.w6(32'h3aeb80b1),
	.w7(32'h3b48ddc6),
	.w8(32'h3beb546e),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bec3bf6),
	.w1(32'h3b87d851),
	.w2(32'hbac0490b),
	.w3(32'h3c7fd625),
	.w4(32'hbb4c85fc),
	.w5(32'hbc133c65),
	.w6(32'h3b1f361a),
	.w7(32'h38122fd3),
	.w8(32'hbc04f1e4),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94e1da4),
	.w1(32'h39e53b1b),
	.w2(32'h3c0434f8),
	.w3(32'h3ba26faa),
	.w4(32'h3b88f3a3),
	.w5(32'hbbf206f4),
	.w6(32'h39eeaecb),
	.w7(32'hbbdfb29d),
	.w8(32'hbbdfaca1),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b32b599),
	.w1(32'h3c68494c),
	.w2(32'h3c06c769),
	.w3(32'h39eba51d),
	.w4(32'h3b5df267),
	.w5(32'h3c75e05d),
	.w6(32'h3bf0d78e),
	.w7(32'h3ba21ba0),
	.w8(32'h3a466d3e),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b892088),
	.w1(32'h3c008678),
	.w2(32'h3bddeda7),
	.w3(32'hbb3687e2),
	.w4(32'h3bf452e6),
	.w5(32'hbc6cba03),
	.w6(32'h3b3c7317),
	.w7(32'hbb24fcc6),
	.w8(32'h3b870997),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a56a43e),
	.w1(32'h3c40afb8),
	.w2(32'hb957adeb),
	.w3(32'hbc1ab842),
	.w4(32'h3bffbe91),
	.w5(32'hbc20d5eb),
	.w6(32'h3b39308c),
	.w7(32'h3b6ffc20),
	.w8(32'h3a1aaa8a),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba7c911),
	.w1(32'h3c8e6c4e),
	.w2(32'hbadfe443),
	.w3(32'hbb8e3806),
	.w4(32'hbb95f12c),
	.w5(32'hbca35c2f),
	.w6(32'h3b41bfef),
	.w7(32'hbbdf7f62),
	.w8(32'hbb75d019),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad89200),
	.w1(32'hbbd3398b),
	.w2(32'h3a94b327),
	.w3(32'h3b295c39),
	.w4(32'h3a094489),
	.w5(32'hbb1e301f),
	.w6(32'hbc3932f9),
	.w7(32'hbae0b595),
	.w8(32'hbaebc514),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba0fd69),
	.w1(32'h3a69f7a5),
	.w2(32'h3a25430b),
	.w3(32'h3bc37a5b),
	.w4(32'h3ac939bd),
	.w5(32'hbbe24166),
	.w6(32'h3b5bde6d),
	.w7(32'hbb3a638e),
	.w8(32'h3a51e1a3),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6faa6f),
	.w1(32'h3b05c94f),
	.w2(32'hbb9b4d26),
	.w3(32'hbafb53b4),
	.w4(32'hbb77ef27),
	.w5(32'h3b53f498),
	.w6(32'h39b13d30),
	.w7(32'h3a5c5696),
	.w8(32'hbab597e0),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc37bf28),
	.w1(32'hbbd80d78),
	.w2(32'hbb4861f5),
	.w3(32'hbc55ca9c),
	.w4(32'hb9d3f7a0),
	.w5(32'hba59cd99),
	.w6(32'hbc128c7c),
	.w7(32'h3b513319),
	.w8(32'h3a3e2132),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcb6501),
	.w1(32'h3ae50fe4),
	.w2(32'hbc4847c6),
	.w3(32'h3afa5dc6),
	.w4(32'h3d152320),
	.w5(32'hbba39166),
	.w6(32'h3bc4aca5),
	.w7(32'h3bf069e0),
	.w8(32'hbb7b5d2a),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba83504e),
	.w1(32'hb9ebcaab),
	.w2(32'hbbadbce6),
	.w3(32'hbc71d622),
	.w4(32'hbb9d6b39),
	.w5(32'hbbeeeebe),
	.w6(32'hbc7eb39e),
	.w7(32'hbb22ec76),
	.w8(32'h3a02f4de),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb04019c),
	.w1(32'hbbc3289f),
	.w2(32'hbc5cfb08),
	.w3(32'hba186787),
	.w4(32'hbb898270),
	.w5(32'hbbc15cdd),
	.w6(32'hbbdf4bc3),
	.w7(32'h3aee2824),
	.w8(32'h3c14c791),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bec1955),
	.w1(32'h3be9b857),
	.w2(32'h3d18a3f9),
	.w3(32'h3c809451),
	.w4(32'h3c0a15a5),
	.w5(32'h3c4fed4a),
	.w6(32'hbb2595e0),
	.w7(32'hbc51640f),
	.w8(32'hbd37158b),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba084dc0),
	.w1(32'h3c12244b),
	.w2(32'hba083274),
	.w3(32'hbb179145),
	.w4(32'h3c58b6eb),
	.w5(32'hbc079539),
	.w6(32'hbad0cd23),
	.w7(32'h3baeee04),
	.w8(32'hbbaf32e5),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6fa2a7),
	.w1(32'h3c14b1e0),
	.w2(32'hbb438525),
	.w3(32'hbc323bdb),
	.w4(32'h3c2c8b72),
	.w5(32'hbcb176d6),
	.w6(32'hbbced692),
	.w7(32'h3c1e2657),
	.w8(32'hbab2e109),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0e28d6),
	.w1(32'hba06d9bd),
	.w2(32'hbb72aa8f),
	.w3(32'hbbad89da),
	.w4(32'h3b9378b8),
	.w5(32'hb981087c),
	.w6(32'hbaaa04f2),
	.w7(32'hbba1a62d),
	.w8(32'hbba6455c),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0be5ba),
	.w1(32'hbc8aa810),
	.w2(32'hba656207),
	.w3(32'hbc6be964),
	.w4(32'hbcfd266f),
	.w5(32'hb9e93185),
	.w6(32'hbc134859),
	.w7(32'hbcb587bc),
	.w8(32'hbb85d7cc),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c063b96),
	.w1(32'h3bd6dc62),
	.w2(32'h3abe935d),
	.w3(32'h3cee13fd),
	.w4(32'h3c53aee2),
	.w5(32'hb9f5da36),
	.w6(32'h3c624693),
	.w7(32'h3b81c9d0),
	.w8(32'h39aaf7a0),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6c3f95),
	.w1(32'hbcf6eadb),
	.w2(32'h3c68ba85),
	.w3(32'hbc662bec),
	.w4(32'hbc04507f),
	.w5(32'h3dad4c56),
	.w6(32'hbc5b2bca),
	.w7(32'hbca504e5),
	.w8(32'hbade335e),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd14941d),
	.w1(32'hbbd81802),
	.w2(32'hbc472265),
	.w3(32'hbd236ae3),
	.w4(32'h3a6ed683),
	.w5(32'hbc56ed0c),
	.w6(32'h3b6b179a),
	.w7(32'hbc2bbc5d),
	.w8(32'hbc9543b4),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7b718b),
	.w1(32'hbc6bc6ce),
	.w2(32'h3be4b7b7),
	.w3(32'hbc8259a9),
	.w4(32'h39e40c53),
	.w5(32'h3ca0bde5),
	.w6(32'hbc613611),
	.w7(32'hbc488815),
	.w8(32'h3c47e191),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b53788e),
	.w1(32'h3b976c85),
	.w2(32'h3c538f48),
	.w3(32'h3a8316db),
	.w4(32'h3ba168c6),
	.w5(32'h3c86fbaf),
	.w6(32'h3c5db0c0),
	.w7(32'h3c0e7352),
	.w8(32'h3c26c174),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2fb8ae),
	.w1(32'h3b4f277e),
	.w2(32'h3b4de468),
	.w3(32'hbb9f44b4),
	.w4(32'h3b1dd668),
	.w5(32'h3c97dbf1),
	.w6(32'hbbc45519),
	.w7(32'hbb966ccd),
	.w8(32'h3bc6cbce),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9401b02),
	.w1(32'h3bea5b86),
	.w2(32'h3b0bddfd),
	.w3(32'h3c3a48a3),
	.w4(32'h3bd1d73d),
	.w5(32'hba81a0c0),
	.w6(32'hbb930d4d),
	.w7(32'h373c3fba),
	.w8(32'h3ac6d5bd),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb3a3cb),
	.w1(32'hba413a77),
	.w2(32'h3c2b9a98),
	.w3(32'h3c0a6bc8),
	.w4(32'hbb8a863e),
	.w5(32'h3b5f6a6c),
	.w6(32'h3aca0107),
	.w7(32'hbc300897),
	.w8(32'hbc956182),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc56641),
	.w1(32'hbc6d577b),
	.w2(32'hbc556efa),
	.w3(32'h398b2dca),
	.w4(32'hbcacd883),
	.w5(32'hbcacad60),
	.w6(32'hbc37d369),
	.w7(32'hbc80849b),
	.w8(32'hbc067049),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8f4ff4),
	.w1(32'hbcad8a00),
	.w2(32'h3c534b0d),
	.w3(32'h3b1ea2a7),
	.w4(32'hbd32f6b4),
	.w5(32'h3cdb2cd3),
	.w6(32'hbb36d817),
	.w7(32'hbcc6d338),
	.w8(32'h3b9303ae),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb36d5f),
	.w1(32'h3c8a2f54),
	.w2(32'hba61ce09),
	.w3(32'h3d2edbeb),
	.w4(32'h3d257aca),
	.w5(32'hbb924693),
	.w6(32'h3c4f2b4f),
	.w7(32'h3c55151f),
	.w8(32'hbc7b2fa2),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd106ba),
	.w1(32'hbb83e48c),
	.w2(32'hb8e50eca),
	.w3(32'hbd708550),
	.w4(32'hbc4adc59),
	.w5(32'hbc3f1913),
	.w6(32'hbd0d5424),
	.w7(32'hbc1d8966),
	.w8(32'hbaf56f1a),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a96812c),
	.w1(32'h3c368b28),
	.w2(32'hba40c98a),
	.w3(32'h3c4bae13),
	.w4(32'h3b5bddad),
	.w5(32'hbbb94036),
	.w6(32'h3b3bbbe8),
	.w7(32'h3c12b89f),
	.w8(32'h3a96bb3e),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2cdec0),
	.w1(32'hbc2f0588),
	.w2(32'hbc0d1905),
	.w3(32'hbb8c154b),
	.w4(32'hbc0ab19e),
	.w5(32'h3b182ba9),
	.w6(32'h39b95fa9),
	.w7(32'hbadb3efe),
	.w8(32'h3c33cb1a),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0b0e25),
	.w1(32'h3b605063),
	.w2(32'hbc58e955),
	.w3(32'h3b9ea036),
	.w4(32'h3b8ea402),
	.w5(32'hbc20c0d9),
	.w6(32'h3b2e28ca),
	.w7(32'h3bee7ae9),
	.w8(32'h3c0a2011),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa80e64),
	.w1(32'hbc262866),
	.w2(32'hbc3ec571),
	.w3(32'hbc20d56b),
	.w4(32'hb91d7734),
	.w5(32'hbc855a53),
	.w6(32'hbbac4083),
	.w7(32'hbc4468ad),
	.w8(32'hbbe6917a),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9c2be0),
	.w1(32'h3ba6e5ad),
	.w2(32'h3a499251),
	.w3(32'hbb696271),
	.w4(32'hba983b66),
	.w5(32'hbc01a431),
	.w6(32'hbc28f20c),
	.w7(32'h3b32efd9),
	.w8(32'hbbd4cb7d),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be5ca15),
	.w1(32'hbb11f74b),
	.w2(32'hb99df343),
	.w3(32'h3b9481e5),
	.w4(32'hbbc25366),
	.w5(32'h3a990088),
	.w6(32'hbb0a231e),
	.w7(32'hbb20f7bf),
	.w8(32'h3b4c117f),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb485065),
	.w1(32'h3b8d038b),
	.w2(32'hbb0039fc),
	.w3(32'hbb73c1e7),
	.w4(32'h3bd9d8e3),
	.w5(32'hbbd16e91),
	.w6(32'hbae1fd39),
	.w7(32'h3bd1f111),
	.w8(32'h3b14e9fb),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbeaab7),
	.w1(32'hbc1248eb),
	.w2(32'hbc2393e1),
	.w3(32'hbbbe1238),
	.w4(32'hbb89962c),
	.w5(32'hbb817b3d),
	.w6(32'hbba700a3),
	.w7(32'hbba314ff),
	.w8(32'hbc14ea9b),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39193fb9),
	.w1(32'h3ae0f6a9),
	.w2(32'hbb2400c6),
	.w3(32'hbbb1e8be),
	.w4(32'h3c16f70b),
	.w5(32'hbbce5adf),
	.w6(32'hbb34d042),
	.w7(32'h3bb3b470),
	.w8(32'h3bcfd53e),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8a1c21),
	.w1(32'h3c42a3ae),
	.w2(32'h3c5aa952),
	.w3(32'h3b1dcd7d),
	.w4(32'hb947de44),
	.w5(32'hbc8f0ec6),
	.w6(32'hbb88c4e4),
	.w7(32'h3bdce30e),
	.w8(32'hbbf48a0a),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd873b1),
	.w1(32'h3a43bada),
	.w2(32'hbbc0c703),
	.w3(32'h3b9e5b93),
	.w4(32'hba9330d6),
	.w5(32'hbc2c789c),
	.w6(32'hbc48896a),
	.w7(32'hbb032ef0),
	.w8(32'hbbe0a903),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b550a81),
	.w1(32'h3bbe0135),
	.w2(32'h3bb533fb),
	.w3(32'h3c0d6eae),
	.w4(32'h3cfa4e7e),
	.w5(32'h3c8a54bd),
	.w6(32'h3afc30f9),
	.w7(32'hbc1e2a9b),
	.w8(32'hbb5d0919),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe1518e),
	.w1(32'hbbc89264),
	.w2(32'h3ad874d2),
	.w3(32'hbc4d2266),
	.w4(32'hbc209002),
	.w5(32'h3c4c6744),
	.w6(32'h3a6f0ced),
	.w7(32'h3adb2e5a),
	.w8(32'h3c155ef9),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b93f290),
	.w1(32'h3b87ff36),
	.w2(32'h3bba611f),
	.w3(32'h3c0d2038),
	.w4(32'h3bc0684d),
	.w5(32'h3bbe7959),
	.w6(32'h3b181015),
	.w7(32'h3b8935fa),
	.w8(32'hbbcfbf6c),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc20884d),
	.w1(32'hbc9dc2e9),
	.w2(32'hbc265f28),
	.w3(32'hbc907574),
	.w4(32'hbcbaac23),
	.w5(32'hbb479bcd),
	.w6(32'hbc4dadb8),
	.w7(32'hbc8e2405),
	.w8(32'hbbb26724),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b43d683),
	.w1(32'h38ad63a2),
	.w2(32'hbc909377),
	.w3(32'h3cbb3ba7),
	.w4(32'hbc3f81ed),
	.w5(32'hbce95b1f),
	.w6(32'h39a3cd6f),
	.w7(32'h3c9acc77),
	.w8(32'h3c8dafe1),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7b9d54),
	.w1(32'h3be16d31),
	.w2(32'hbbd2e472),
	.w3(32'h3cbe0f0d),
	.w4(32'h3b9564bd),
	.w5(32'hbcf873cf),
	.w6(32'h3c688871),
	.w7(32'h3c16c1ee),
	.w8(32'hba568220),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb40c2d9),
	.w1(32'h3acb6c4b),
	.w2(32'h3b447b4e),
	.w3(32'hbc370dd2),
	.w4(32'h3c549cf1),
	.w5(32'hba3fd3f5),
	.w6(32'hbc1a8a33),
	.w7(32'h3b4a3400),
	.w8(32'h3a96d5e9),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba58a8c8),
	.w1(32'h3bd424ad),
	.w2(32'h3ba0d510),
	.w3(32'hbaab82bc),
	.w4(32'h3bee32b3),
	.w5(32'hbc46115a),
	.w6(32'hbc0a77c8),
	.w7(32'h3c2ad299),
	.w8(32'hbb96b7ea),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b935eb7),
	.w1(32'hbc1ebf33),
	.w2(32'hbbdeb0a9),
	.w3(32'h3c7a65c5),
	.w4(32'hbc3c4761),
	.w5(32'hbba4141c),
	.w6(32'h3c03b330),
	.w7(32'hbbfd9b08),
	.w8(32'hbbad3d91),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb795407),
	.w1(32'hbc0beeed),
	.w2(32'h3b140be6),
	.w3(32'hbc18a8d1),
	.w4(32'hbb47ba14),
	.w5(32'h3b1cccf6),
	.w6(32'h3b07fddd),
	.w7(32'hbba6e154),
	.w8(32'hbaa29aee),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb57c515),
	.w1(32'hba98139e),
	.w2(32'h3b627329),
	.w3(32'hbb66f1f1),
	.w4(32'h3b04e9eb),
	.w5(32'hbbd1ba6e),
	.w6(32'h3b2aca36),
	.w7(32'hbb3baa53),
	.w8(32'hbbafc517),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1b13e3),
	.w1(32'hba4a3fac),
	.w2(32'hbb84742d),
	.w3(32'h3c3163a0),
	.w4(32'hba1e7c27),
	.w5(32'h3b992016),
	.w6(32'h3b16dbb5),
	.w7(32'h3aa085b4),
	.w8(32'h3be3a978),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0ad120),
	.w1(32'h3bf7ddb0),
	.w2(32'h3aac2a23),
	.w3(32'hbb4bc3cf),
	.w4(32'hbb6c3dde),
	.w5(32'h39df7d4e),
	.w6(32'h3b8dd988),
	.w7(32'h3b35010e),
	.w8(32'hbb820710),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7bd0d5),
	.w1(32'hb81404e5),
	.w2(32'hbc12d25a),
	.w3(32'h3abd9388),
	.w4(32'hbac03c9a),
	.w5(32'h3bdce48f),
	.w6(32'hbbaaf58d),
	.w7(32'hbb9c6b83),
	.w8(32'hbac2b9f4),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf371ef),
	.w1(32'hba3100f3),
	.w2(32'h3b569d07),
	.w3(32'h3b216861),
	.w4(32'hbaa60f68),
	.w5(32'hb99babbc),
	.w6(32'h3be596b2),
	.w7(32'h3accdc26),
	.w8(32'h3a997976),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd7782b),
	.w1(32'h3afee9b2),
	.w2(32'h3bc6505f),
	.w3(32'h3ab68f21),
	.w4(32'hbbcfe97d),
	.w5(32'h3cb1ff64),
	.w6(32'h3b7320fb),
	.w7(32'hbc4c2c0e),
	.w8(32'hbb0977a4),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b811295),
	.w1(32'hbb5298f5),
	.w2(32'hbb7568a4),
	.w3(32'hba75b8cc),
	.w4(32'hbbd910d5),
	.w5(32'h3a98e267),
	.w6(32'h3b2e6148),
	.w7(32'hba2154e9),
	.w8(32'h39f32a2b),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5349a7),
	.w1(32'hbb6736a5),
	.w2(32'h3a2d77fe),
	.w3(32'h3b457eb1),
	.w4(32'h3b852632),
	.w5(32'hba9ebd48),
	.w6(32'h3a012023),
	.w7(32'h3b52f4e6),
	.w8(32'hbb599bba),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2fd15b),
	.w1(32'h3b9aacb4),
	.w2(32'hb991d910),
	.w3(32'hbbea480a),
	.w4(32'h3b3e241d),
	.w5(32'h3a1b2249),
	.w6(32'hbb7c2a93),
	.w7(32'h3c0f4ecc),
	.w8(32'h3c0e7010),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacf8caa),
	.w1(32'h3aa72e7a),
	.w2(32'hbacc81e7),
	.w3(32'hb9df29cf),
	.w4(32'h3a5c931c),
	.w5(32'h3bd1c3a0),
	.w6(32'h3c21f775),
	.w7(32'hbb1a5c98),
	.w8(32'h39a75c12),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2ae291),
	.w1(32'h39ce12b3),
	.w2(32'h3c0b8c92),
	.w3(32'hbc051e46),
	.w4(32'h3baddd36),
	.w5(32'h3b91cbae),
	.w6(32'hb9c27624),
	.w7(32'h3befcc22),
	.w8(32'h3b7ca04b),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b80c2c4),
	.w1(32'h3c0fc83b),
	.w2(32'h3a97045d),
	.w3(32'hb9f05071),
	.w4(32'h3ba76967),
	.w5(32'h3b1368be),
	.w6(32'hbae29fcf),
	.w7(32'h3a6cfa1f),
	.w8(32'h3bd57120),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7c661b),
	.w1(32'h3b2daac1),
	.w2(32'hbb50b8dd),
	.w3(32'h3c209b9d),
	.w4(32'hbbca92c3),
	.w5(32'h3b8addfc),
	.w6(32'h3c1c2506),
	.w7(32'h3a9c54e1),
	.w8(32'h383700b5),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390a6f61),
	.w1(32'hbc043e81),
	.w2(32'h3b68626a),
	.w3(32'h3969966f),
	.w4(32'hbbd5056f),
	.w5(32'h3c893d47),
	.w6(32'h3a125dbe),
	.w7(32'h3bb8a873),
	.w8(32'h3a9988e3),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c439b06),
	.w1(32'hbb2eb64c),
	.w2(32'hbbb718b1),
	.w3(32'h3c5f3b1e),
	.w4(32'h39a64362),
	.w5(32'hbc365b5b),
	.w6(32'hbba09d6a),
	.w7(32'hbb2c98b1),
	.w8(32'h3b44aea6),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae1ac83),
	.w1(32'h3a999803),
	.w2(32'h3b80062a),
	.w3(32'hbbeca2ff),
	.w4(32'hbb188eaa),
	.w5(32'h3b275379),
	.w6(32'hbc151ffe),
	.w7(32'h3942dae5),
	.w8(32'h3952c9fa),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acadc82),
	.w1(32'hbb7355bd),
	.w2(32'hbba1937e),
	.w3(32'hbb201254),
	.w4(32'hbb4673a9),
	.w5(32'hbb350cbf),
	.w6(32'hbc5a7bda),
	.w7(32'hbb943046),
	.w8(32'hbbed1d1e),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb996202),
	.w1(32'h3c3befad),
	.w2(32'h3c1da480),
	.w3(32'hbc125c29),
	.w4(32'h3cbef78c),
	.w5(32'h3c1b59ee),
	.w6(32'h3bd3ddf6),
	.w7(32'h3b8ab134),
	.w8(32'h3c866836),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3825dc),
	.w1(32'hb9ed1376),
	.w2(32'hbb508f30),
	.w3(32'hbb3761c9),
	.w4(32'hbab9879e),
	.w5(32'hbc1a78b6),
	.w6(32'h3c64a398),
	.w7(32'hbb1a2b12),
	.w8(32'hbbcc40f3),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b5872),
	.w1(32'hbb2764cf),
	.w2(32'h3b9c3974),
	.w3(32'hbc46d7ad),
	.w4(32'hbaa25aa3),
	.w5(32'h3c400b5e),
	.w6(32'h3b3a313e),
	.w7(32'hbb4e9181),
	.w8(32'hbaab4430),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aca0540),
	.w1(32'h3bf2b701),
	.w2(32'h3b89b504),
	.w3(32'h3be4fdb7),
	.w4(32'h3b07cb75),
	.w5(32'hbb6ebafd),
	.w6(32'h392a32ed),
	.w7(32'h3c1c7924),
	.w8(32'hbbcf9933),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a25445a),
	.w1(32'h3b0b58c1),
	.w2(32'h3baf458f),
	.w3(32'hbb280164),
	.w4(32'h3b543f62),
	.w5(32'h3a4bcc30),
	.w6(32'hbaaeb3a6),
	.w7(32'h3bda091a),
	.w8(32'h3a45ba91),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h378d3902),
	.w1(32'hbad80782),
	.w2(32'h3b450b07),
	.w3(32'h3b9d9035),
	.w4(32'h3b9f7e86),
	.w5(32'hbbfccd4c),
	.w6(32'h3a437948),
	.w7(32'h3b996c01),
	.w8(32'h3bcc1d70),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf0ab82),
	.w1(32'h3b01a792),
	.w2(32'h3ada9957),
	.w3(32'hbbd9d25e),
	.w4(32'h3b550424),
	.w5(32'hbb640685),
	.w6(32'hbb984519),
	.w7(32'hbbe8d77e),
	.w8(32'hbb22e399),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7de50f),
	.w1(32'hbb5e7ba4),
	.w2(32'h3b832dc1),
	.w3(32'hbb7e39db),
	.w4(32'hbbba1e6a),
	.w5(32'h3c7aa3ea),
	.w6(32'hbb62bd26),
	.w7(32'h3bc9ba8d),
	.w8(32'h3bea28aa),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2342d1),
	.w1(32'h3c8b2bdb),
	.w2(32'h3abf83b5),
	.w3(32'h3afc418e),
	.w4(32'h3c81ef91),
	.w5(32'h3c1e701f),
	.w6(32'h3a061c5a),
	.w7(32'h3ba5649b),
	.w8(32'h3bb8b2b2),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afd383e),
	.w1(32'h3b1e193c),
	.w2(32'h3aa51a61),
	.w3(32'hbb8057d3),
	.w4(32'h3ca948b4),
	.w5(32'hbc06bcf2),
	.w6(32'h3c1d2f77),
	.w7(32'h3b6608be),
	.w8(32'h3c29534f),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bad47f5),
	.w1(32'h3bede56e),
	.w2(32'h3b145505),
	.w3(32'hb9584ed0),
	.w4(32'h3c0d4630),
	.w5(32'h3ce34986),
	.w6(32'h3bf1da3a),
	.w7(32'hbc13a7ed),
	.w8(32'hbb8c6243),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396ce7c6),
	.w1(32'hbbe649ff),
	.w2(32'hbba9e30f),
	.w3(32'h3c390e07),
	.w4(32'hbb6d71cc),
	.w5(32'hbbac858c),
	.w6(32'h3bcf73e3),
	.w7(32'hba930ddd),
	.w8(32'hbafa56dd),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba839c08),
	.w1(32'h3b07ad2a),
	.w2(32'h3ac94cb3),
	.w3(32'hbbdb98cc),
	.w4(32'hbc1981e9),
	.w5(32'h3bee6526),
	.w6(32'hba8ac015),
	.w7(32'h3a6880bd),
	.w8(32'hbb96180f),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8eaffe),
	.w1(32'hbc120a4e),
	.w2(32'hbaf3fbc5),
	.w3(32'h3c180351),
	.w4(32'hbb788b85),
	.w5(32'h3b61cf3f),
	.w6(32'hb9a55866),
	.w7(32'hbbe272be),
	.w8(32'h39b048b2),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a67dabc),
	.w1(32'h3ba6baee),
	.w2(32'h3af49472),
	.w3(32'hbaacf6f6),
	.w4(32'hba94a501),
	.w5(32'h3bc854e5),
	.w6(32'hbb1309b0),
	.w7(32'hbac3850d),
	.w8(32'h3a56358e),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf22799),
	.w1(32'hbb13a10f),
	.w2(32'hba99e1e9),
	.w3(32'h38c0ee68),
	.w4(32'h38128eb3),
	.w5(32'h3b013c9c),
	.w6(32'h3ba91b60),
	.w7(32'hbb72dd6e),
	.w8(32'hbb264b44),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbc67a0),
	.w1(32'hbb255480),
	.w2(32'hbb9757ab),
	.w3(32'hbbf3aa13),
	.w4(32'hba9584a8),
	.w5(32'hbb44d3ba),
	.w6(32'hbb644048),
	.w7(32'hba5b0c28),
	.w8(32'h3aceeee5),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b246ace),
	.w1(32'hbb4fbc9d),
	.w2(32'h3a868a1d),
	.w3(32'h3af03b89),
	.w4(32'h3b12b7ad),
	.w5(32'h3c007503),
	.w6(32'h3ac035e3),
	.w7(32'hbb76af3d),
	.w8(32'hbb803917),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3ca0c5),
	.w1(32'h3b4f6f16),
	.w2(32'hbbaf495e),
	.w3(32'hba8e30df),
	.w4(32'hbb3d513f),
	.w5(32'hba3a8345),
	.w6(32'hbb8f1a2e),
	.w7(32'h3b949356),
	.w8(32'h3b2d04cf),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa32740),
	.w1(32'h3bcebc9a),
	.w2(32'h3c1c421b),
	.w3(32'hbb9b5d1e),
	.w4(32'h3bf67014),
	.w5(32'h3c0d352b),
	.w6(32'hb96c91d2),
	.w7(32'hbbc21813),
	.w8(32'h3be58e75),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfcacb5),
	.w1(32'h3b0a5506),
	.w2(32'hbb0bfe71),
	.w3(32'hb8a50e7b),
	.w4(32'h3bcb64b7),
	.w5(32'hbba73c7b),
	.w6(32'h3c141b8a),
	.w7(32'h3be16032),
	.w8(32'hba9b97ff),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2782dd),
	.w1(32'h3b047b1f),
	.w2(32'h3c05ee73),
	.w3(32'hbb2c5736),
	.w4(32'h3ce2e7d2),
	.w5(32'h3c45dbb8),
	.w6(32'hbbfc5d15),
	.w7(32'h3c039709),
	.w8(32'hbaa6a252),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b892467),
	.w1(32'h3c33bb17),
	.w2(32'h3c6060b3),
	.w3(32'hbb5bf52b),
	.w4(32'h3c525291),
	.w5(32'h3b5ba4cd),
	.w6(32'h3af92cae),
	.w7(32'h3b9943da),
	.w8(32'h3c2505e0),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b431649),
	.w1(32'h3b69d424),
	.w2(32'h3c0780b9),
	.w3(32'h3bcfd383),
	.w4(32'hbc0bed4e),
	.w5(32'h3c66d5b7),
	.w6(32'h3bb75121),
	.w7(32'h3b5df269),
	.w8(32'h3be4721d),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbd8875),
	.w1(32'hbb6fd0e2),
	.w2(32'h3b541cfb),
	.w3(32'h3b8e2934),
	.w4(32'hbbac2c93),
	.w5(32'h3b7f4e43),
	.w6(32'h3c2ec4f6),
	.w7(32'h3bcdfcfa),
	.w8(32'hbaae9520),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b04f521),
	.w1(32'h3a27aaf7),
	.w2(32'h3c04898b),
	.w3(32'hba3bb031),
	.w4(32'h3ba532a4),
	.w5(32'h3b30646a),
	.w6(32'h3a848fc3),
	.w7(32'h3c1fbb4f),
	.w8(32'h3bb45b9b),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c155144),
	.w1(32'hbbc9e89d),
	.w2(32'hbb08f5d4),
	.w3(32'h3c837db0),
	.w4(32'hbbfa6078),
	.w5(32'h3b9e88c3),
	.w6(32'h3bc64dc8),
	.w7(32'hbb605b55),
	.w8(32'h3ad0c059),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb78b4b4),
	.w1(32'h3b272374),
	.w2(32'h3c17d423),
	.w3(32'h3ac32035),
	.w4(32'h3b178d36),
	.w5(32'h3bc7cd07),
	.w6(32'h3b9d48aa),
	.w7(32'h3b875c9b),
	.w8(32'h3af9a3fe),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd52617),
	.w1(32'hbae8a219),
	.w2(32'h3b7ddda8),
	.w3(32'h3c83691a),
	.w4(32'h3b5e9ac2),
	.w5(32'h3ad26d1b),
	.w6(32'h3c036707),
	.w7(32'h3a886b46),
	.w8(32'h3bc56759),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc1f96e),
	.w1(32'hbba72bce),
	.w2(32'hbb8b6f24),
	.w3(32'hbba1acca),
	.w4(32'hbc157f48),
	.w5(32'hbab0c90b),
	.w6(32'hba90c8f8),
	.w7(32'hbc3a5596),
	.w8(32'hbc0ffa5d),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af57754),
	.w1(32'hbbf4b7c1),
	.w2(32'hbb051954),
	.w3(32'hbb7f4000),
	.w4(32'hbb865534),
	.w5(32'hbb9e9a80),
	.w6(32'hba869276),
	.w7(32'hbba9ae12),
	.w8(32'h3b150661),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae72083),
	.w1(32'hba982d89),
	.w2(32'hb98a4e75),
	.w3(32'hbba3c56f),
	.w4(32'hbb4cf3ac),
	.w5(32'h3b1cfebf),
	.w6(32'h3a48560e),
	.w7(32'hbb2bf048),
	.w8(32'hbb9cd8a8),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6a5eb5),
	.w1(32'h3ae519b0),
	.w2(32'h3be3f46f),
	.w3(32'h390d0310),
	.w4(32'h3b988d9c),
	.w5(32'hbb88081d),
	.w6(32'h3b493927),
	.w7(32'hbb17c680),
	.w8(32'hbb4fc173),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbae625),
	.w1(32'hbbec819f),
	.w2(32'h3a6fdf96),
	.w3(32'h3ae97350),
	.w4(32'hbc0ef012),
	.w5(32'h3c2f3bf3),
	.w6(32'h3b2b5fd4),
	.w7(32'hbb2202cf),
	.w8(32'h3ab0bb71),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a684f0d),
	.w1(32'hbaa042b5),
	.w2(32'hbbe9cbe9),
	.w3(32'h3c093192),
	.w4(32'hbba3a2ee),
	.w5(32'h3b8f5e30),
	.w6(32'h3a344f68),
	.w7(32'h3bced338),
	.w8(32'hba11a54f),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc071e4d),
	.w1(32'hbc0884b9),
	.w2(32'h3802f272),
	.w3(32'h3aef8b93),
	.w4(32'hbc0799dc),
	.w5(32'h3be1e263),
	.w6(32'h3a1a29dc),
	.w7(32'hbc305114),
	.w8(32'hbb99f830),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb28f102),
	.w1(32'hbb6a580f),
	.w2(32'hbac779a2),
	.w3(32'h3b38ff58),
	.w4(32'hbbe5ddc5),
	.w5(32'hb9d07fb1),
	.w6(32'hba8a08b6),
	.w7(32'hbb3d246c),
	.w8(32'hbc0a6056),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a101d0d),
	.w1(32'hba3f7ca4),
	.w2(32'hba5e461e),
	.w3(32'h3aa016db),
	.w4(32'hbb334ec0),
	.w5(32'hbc475777),
	.w6(32'hbc1a862b),
	.w7(32'hbb1ef8c7),
	.w8(32'h3a86b3ff),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdf55db),
	.w1(32'h3a87bbbc),
	.w2(32'hbb5a7989),
	.w3(32'h3a0face7),
	.w4(32'hbbf47828),
	.w5(32'h3c2ee22b),
	.w6(32'hbb940426),
	.w7(32'hbaf2f145),
	.w8(32'h3c58c5a3),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad98211),
	.w1(32'hb9bc0a23),
	.w2(32'hbaaf6277),
	.w3(32'h3c1510b9),
	.w4(32'hbbb4e249),
	.w5(32'hbc1881a3),
	.w6(32'h3ab6b0f9),
	.w7(32'h389d2197),
	.w8(32'h3ae70c99),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aac1fa8),
	.w1(32'hbaa8e33d),
	.w2(32'h3b9c8149),
	.w3(32'hbba48e64),
	.w4(32'hbb5d47aa),
	.w5(32'h3bdc0165),
	.w6(32'h39861dc5),
	.w7(32'hba5ad64b),
	.w8(32'h3b7ae3a3),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd4666b),
	.w1(32'h3abd25f9),
	.w2(32'hbb6c14e6),
	.w3(32'h3ba8028d),
	.w4(32'h3bcd853a),
	.w5(32'hbad370dd),
	.w6(32'h3b91dd4e),
	.w7(32'h3afe5416),
	.w8(32'hbab76f4a),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac6b13d),
	.w1(32'hbb7a91e7),
	.w2(32'h3a4870e7),
	.w3(32'hbb5ead91),
	.w4(32'hbaf5259f),
	.w5(32'h3b70b3d2),
	.w6(32'h3a46c8cd),
	.w7(32'hbbc74e07),
	.w8(32'hbb0900b7),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88b38d7),
	.w1(32'h3b10771b),
	.w2(32'h3a08115c),
	.w3(32'h3c06c3bc),
	.w4(32'h39898f85),
	.w5(32'hb9f6d772),
	.w6(32'h3b82b16f),
	.w7(32'h3b9a7994),
	.w8(32'h3b223eae),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb59b4f7a),
	.w1(32'h3b5402d7),
	.w2(32'h3b9313d0),
	.w3(32'h3afd256e),
	.w4(32'hbc4c8b42),
	.w5(32'h3c79c58a),
	.w6(32'h3bb92e7a),
	.w7(32'h3a8b1e18),
	.w8(32'h3b543986),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaf8b90),
	.w1(32'h3b6446fb),
	.w2(32'hbb2698c3),
	.w3(32'h3c6eb62a),
	.w4(32'hbb8908b1),
	.w5(32'hb8d4abf4),
	.w6(32'h3a7a19e3),
	.w7(32'hbbaf3cbd),
	.w8(32'hbb170029),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5c6f89),
	.w1(32'h3a910c99),
	.w2(32'h3bf3f691),
	.w3(32'hbbdf1b95),
	.w4(32'h3c1fd4b7),
	.w5(32'h39cb8a07),
	.w6(32'hbb85935d),
	.w7(32'h3bcd8475),
	.w8(32'h386b4e8f),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abc8712),
	.w1(32'h3b05b16e),
	.w2(32'h3b20c679),
	.w3(32'hbb6e4150),
	.w4(32'h3aa652c6),
	.w5(32'h3b4546b7),
	.w6(32'hbb158aaf),
	.w7(32'h3b7ef3e6),
	.w8(32'h3bba4cc2),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc7d07d),
	.w1(32'h3ad70d69),
	.w2(32'h3c1e46fb),
	.w3(32'h3b290c63),
	.w4(32'h3b5f5e6a),
	.w5(32'h3b2babc0),
	.w6(32'h3bc0e690),
	.w7(32'h3b16399b),
	.w8(32'hb98143d5),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be10c9a),
	.w1(32'hb9325109),
	.w2(32'h3b00da57),
	.w3(32'hbb3d5743),
	.w4(32'h3b1eb89e),
	.w5(32'h3c36e0ce),
	.w6(32'hbb9b04c7),
	.w7(32'hbad3175c),
	.w8(32'h3ad815d6),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d24f8),
	.w1(32'hba2fcaf1),
	.w2(32'hbba44f51),
	.w3(32'hbb4b53b9),
	.w4(32'hb9273b12),
	.w5(32'h3a8a0a53),
	.w6(32'h37d8caca),
	.w7(32'h38916429),
	.w8(32'h3b0aac4a),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcd5223),
	.w1(32'hbbaafb31),
	.w2(32'h3bccc655),
	.w3(32'hbbc2575f),
	.w4(32'hbbbf1cc1),
	.w5(32'h3c8e9cf5),
	.w6(32'hbb8a6be9),
	.w7(32'h39cf32f4),
	.w8(32'h3a964e35),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a895bf),
	.w1(32'h3b449f4c),
	.w2(32'hbbc5a87b),
	.w3(32'hbae52bf1),
	.w4(32'hb8cc1ef6),
	.w5(32'hbbe52634),
	.w6(32'hbbad7667),
	.w7(32'hbb821f44),
	.w8(32'h3b20f1f3),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7996ec),
	.w1(32'h3a0b5f65),
	.w2(32'h3bbf38ed),
	.w3(32'h3b4296ab),
	.w4(32'hbc2b73b8),
	.w5(32'h3cc9353e),
	.w6(32'h3b20dbe2),
	.w7(32'hbbf0d5a2),
	.w8(32'h3b4f8352),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c08c58a),
	.w1(32'hbc290c55),
	.w2(32'hbc6003c9),
	.w3(32'h3c34d7af),
	.w4(32'hbc2088b3),
	.w5(32'h3bb9216b),
	.w6(32'h3bf46383),
	.w7(32'hbc04020f),
	.w8(32'hbb4c8e77),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8603e1),
	.w1(32'hbac54a1c),
	.w2(32'h3c2495c0),
	.w3(32'h3ac4aa30),
	.w4(32'hbbd92fab),
	.w5(32'hbb4ef30d),
	.w6(32'h3b3df826),
	.w7(32'hbbb47e69),
	.w8(32'hbb01b187),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfb03e5),
	.w1(32'hba26d12f),
	.w2(32'h3b77a010),
	.w3(32'hba32e035),
	.w4(32'hbba9b462),
	.w5(32'hbc03100a),
	.w6(32'hbacf7693),
	.w7(32'hb9e9f935),
	.w8(32'h38e3ea2b),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c034d33),
	.w1(32'hbb1004c9),
	.w2(32'hb853ba81),
	.w3(32'h3add9cbb),
	.w4(32'hbc28d27b),
	.w5(32'h3bf94722),
	.w6(32'hbafdd261),
	.w7(32'hbb4a80a5),
	.w8(32'hbadbe0b4),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad1b7bf),
	.w1(32'h3c42f3fa),
	.w2(32'h3c0ca165),
	.w3(32'hbace655b),
	.w4(32'hbbba0845),
	.w5(32'h3c921a5b),
	.w6(32'h3b8cb5b2),
	.w7(32'h3b15ca7b),
	.w8(32'hbc673994),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2a7fa3),
	.w1(32'h3a6cb847),
	.w2(32'h3c42aa4f),
	.w3(32'h3c3e2929),
	.w4(32'hbb9ee390),
	.w5(32'h3c568623),
	.w6(32'h3a144d51),
	.w7(32'h3ac4f152),
	.w8(32'h3b03bd35),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5c9626),
	.w1(32'h3c259f74),
	.w2(32'h3c04734c),
	.w3(32'h3639b116),
	.w4(32'hbbc6923d),
	.w5(32'h3cd08c8b),
	.w6(32'hbb70aa57),
	.w7(32'h3ac5af9a),
	.w8(32'h3b4d17c3),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c743943),
	.w1(32'h390cb945),
	.w2(32'h3b990385),
	.w3(32'h3ccf74fd),
	.w4(32'h3b4d8f89),
	.w5(32'hbb999ca6),
	.w6(32'h3ba26873),
	.w7(32'hbb50e99b),
	.w8(32'hb72f204b),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb036d4d),
	.w1(32'h3b8ced0b),
	.w2(32'h3bd9ae14),
	.w3(32'hbaded4c2),
	.w4(32'hbb926daa),
	.w5(32'hbb17489d),
	.w6(32'h3ab5bb69),
	.w7(32'hba2c45e0),
	.w8(32'hbaf7fd12),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab40f5d),
	.w1(32'h3b540330),
	.w2(32'h3ae04019),
	.w3(32'hba43a895),
	.w4(32'h3be9d44f),
	.w5(32'hbbeab209),
	.w6(32'hba01e285),
	.w7(32'h3bcb3680),
	.w8(32'hbbe534ce),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b27cee1),
	.w1(32'h3c19ac08),
	.w2(32'h3c657b77),
	.w3(32'h3c697c3a),
	.w4(32'hba2f8913),
	.w5(32'h3bb07d93),
	.w6(32'h3bfc148c),
	.w7(32'h396c682f),
	.w8(32'h3be17ac3),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c969fc2),
	.w1(32'h3bee368d),
	.w2(32'hbb0c7b08),
	.w3(32'h3cec3195),
	.w4(32'hbc37c7fb),
	.w5(32'h3b4edd6f),
	.w6(32'h3c823e5b),
	.w7(32'hbc12f92e),
	.w8(32'h3a461bbf),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b31c4e6),
	.w1(32'h3b664849),
	.w2(32'h3bb06af1),
	.w3(32'h3b931c6d),
	.w4(32'h3c0bc06b),
	.w5(32'hbbace9c6),
	.w6(32'hb9df5e2e),
	.w7(32'hbb4d081c),
	.w8(32'hba9f6d48),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb627c7b),
	.w1(32'h3c2a6d4f),
	.w2(32'hbb437f21),
	.w3(32'hbbb84180),
	.w4(32'h3b0e9c9f),
	.w5(32'hbc15e827),
	.w6(32'h3a556343),
	.w7(32'hbc0a9a0b),
	.w8(32'hbbf51cfa),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4c505b),
	.w1(32'h3bbefc8c),
	.w2(32'hba0cc348),
	.w3(32'hbc079010),
	.w4(32'h3bfb146b),
	.w5(32'h3b975c28),
	.w6(32'h3be46341),
	.w7(32'h3b997077),
	.w8(32'h3b7ca257),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc724582),
	.w1(32'h3997ebe1),
	.w2(32'h3c03499b),
	.w3(32'hbc6df8d5),
	.w4(32'hbbc66448),
	.w5(32'h3b400735),
	.w6(32'hbb332123),
	.w7(32'hbc07fcbc),
	.w8(32'hbbce1146),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b099162),
	.w1(32'h3b914a4b),
	.w2(32'h3ac3b7e7),
	.w3(32'hbb591c5e),
	.w4(32'h3c2a7257),
	.w5(32'h3bd36f02),
	.w6(32'hbc08ab8c),
	.w7(32'h3b7e7c3c),
	.w8(32'h3ba48160),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb96416),
	.w1(32'hb80200e1),
	.w2(32'hbafd5981),
	.w3(32'h3b704444),
	.w4(32'h3c517ff9),
	.w5(32'hbb71862d),
	.w6(32'h3b691f21),
	.w7(32'h3bfeda87),
	.w8(32'h3c85b824),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba609121),
	.w1(32'h3c33645f),
	.w2(32'h3c3f1f41),
	.w3(32'hbbd4b582),
	.w4(32'h3c891b69),
	.w5(32'h3c45645a),
	.w6(32'h3c00b738),
	.w7(32'h3b098b4a),
	.w8(32'h3bd4b841),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa2a1b7),
	.w1(32'h3b4012b1),
	.w2(32'h3b48b156),
	.w3(32'hba30b1ac),
	.w4(32'h3b466ad2),
	.w5(32'hbbfa8295),
	.w6(32'h3c4b647c),
	.w7(32'hbafc9d00),
	.w8(32'hbb168250),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb368992),
	.w1(32'hbb0475e5),
	.w2(32'hbbd44e68),
	.w3(32'hbb8eeca8),
	.w4(32'hbb4ca69e),
	.w5(32'hbbecd8c2),
	.w6(32'h39fc2f9e),
	.w7(32'hba27ce45),
	.w8(32'hbb990431),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba24b453),
	.w1(32'hba531921),
	.w2(32'hbbc40f92),
	.w3(32'hba6a825b),
	.w4(32'h3a8051a8),
	.w5(32'h3c0dc73a),
	.w6(32'h3975fc72),
	.w7(32'h3b3b5f24),
	.w8(32'hbb1a03e6),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2c9ccd),
	.w1(32'hbb18637c),
	.w2(32'hbc006e25),
	.w3(32'hbae382cf),
	.w4(32'h39f14b14),
	.w5(32'h3976caed),
	.w6(32'hb836ec41),
	.w7(32'hba1c26a5),
	.w8(32'hbbc80f05),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9ce167),
	.w1(32'hbabe27ac),
	.w2(32'hba42ec64),
	.w3(32'hbaf518c3),
	.w4(32'h3b2218e3),
	.w5(32'hbc2e1946),
	.w6(32'hbad3bb22),
	.w7(32'hbb935fa7),
	.w8(32'hbaf074cc),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e82965),
	.w1(32'h3b74e04e),
	.w2(32'h3bb53867),
	.w3(32'hbbd2dd64),
	.w4(32'hbb631304),
	.w5(32'hbb1d51df),
	.w6(32'hbbe5ca08),
	.w7(32'h3a1cf85a),
	.w8(32'h3baa8947),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2ac48e),
	.w1(32'hbbc10888),
	.w2(32'hba4e5e1b),
	.w3(32'h3be5c7e6),
	.w4(32'hbb4965cf),
	.w5(32'h3c2926f0),
	.w6(32'h3bc1aca0),
	.w7(32'hbb8fa0a2),
	.w8(32'hbb2208c2),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5495ba),
	.w1(32'hbb9872a3),
	.w2(32'h3bea8bf6),
	.w3(32'h3b3bd157),
	.w4(32'hbbfebab2),
	.w5(32'h3c962299),
	.w6(32'h3b83c55f),
	.w7(32'hbb47ae1e),
	.w8(32'h3adc7986),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafa89f1),
	.w1(32'h3ac513a5),
	.w2(32'h3b46a60f),
	.w3(32'hba885997),
	.w4(32'h3b88953d),
	.w5(32'h3b8960cb),
	.w6(32'hbbb11cd7),
	.w7(32'h3baae4fb),
	.w8(32'hba4bf386),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c02adb5),
	.w1(32'h39da48a3),
	.w2(32'h3b75233a),
	.w3(32'h3be0cd97),
	.w4(32'h3ac05302),
	.w5(32'hbb3daa42),
	.w6(32'h3bfe999a),
	.w7(32'hbaad0fbb),
	.w8(32'h3be8addc),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b207a63),
	.w1(32'hbbcf15d5),
	.w2(32'h3b6c489c),
	.w3(32'h3a28528a),
	.w4(32'hbc3f7aa6),
	.w5(32'h3b758244),
	.w6(32'h3ba1167a),
	.w7(32'hbbfd525e),
	.w8(32'hbbbfc06e),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3b0091),
	.w1(32'hbb858fe9),
	.w2(32'hbb9cac2c),
	.w3(32'h3b055367),
	.w4(32'hbb281a41),
	.w5(32'h3c06f678),
	.w6(32'h3b9d2f22),
	.w7(32'hbbe440fb),
	.w8(32'h35987b2f),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc4abd6),
	.w1(32'hbbb442ad),
	.w2(32'h3b2683e6),
	.w3(32'hbb640fca),
	.w4(32'h399cd348),
	.w5(32'h3c46a101),
	.w6(32'hbb591dac),
	.w7(32'h3c21e615),
	.w8(32'h38f475ae),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2d5ec4),
	.w1(32'hb8e4f9b4),
	.w2(32'hbb3d4541),
	.w3(32'h3b8278de),
	.w4(32'h3bfc7742),
	.w5(32'hbc18027a),
	.w6(32'hbc25bdef),
	.w7(32'hb94b071d),
	.w8(32'hbb44fdcc),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0754c3),
	.w1(32'h3b627c3e),
	.w2(32'h3b806001),
	.w3(32'hbc274ded),
	.w4(32'h3add1ff0),
	.w5(32'hbbc43d0f),
	.w6(32'hbc047824),
	.w7(32'h3b49780d),
	.w8(32'hba522265),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9d434f),
	.w1(32'h3a1568d8),
	.w2(32'h3bbdb5c5),
	.w3(32'h3b090465),
	.w4(32'h3c1757d2),
	.w5(32'hbaaac992),
	.w6(32'h39e6e2d5),
	.w7(32'h3b291b99),
	.w8(32'hbb592f81),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbe2560),
	.w1(32'hba1a120d),
	.w2(32'hbb974259),
	.w3(32'h3b004363),
	.w4(32'hbb88421f),
	.w5(32'hbc64eeb0),
	.w6(32'h3b4cc7f1),
	.w7(32'hbb1dddff),
	.w8(32'hbbfdac9c),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae1e3fb),
	.w1(32'h3a83a63d),
	.w2(32'h3a10c438),
	.w3(32'h3ac00499),
	.w4(32'hbb7f4a7a),
	.w5(32'h3c0d4586),
	.w6(32'h3bb6a94d),
	.w7(32'h3b122cfe),
	.w8(32'h395a925e),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf77b09),
	.w1(32'h3b84ddf5),
	.w2(32'h3a9aef60),
	.w3(32'h3b6e8cb4),
	.w4(32'h396c1374),
	.w5(32'hbac62525),
	.w6(32'h3bbf2e8e),
	.w7(32'hbab54582),
	.w8(32'h3bd4a826),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2ba8af),
	.w1(32'h3aa840e0),
	.w2(32'h3b898c70),
	.w3(32'h3b929a4c),
	.w4(32'hb9148737),
	.w5(32'hbba09541),
	.w6(32'h3bdd5693),
	.w7(32'h3bf6cd13),
	.w8(32'h3b1dc48d),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5cafae),
	.w1(32'hbbc3e456),
	.w2(32'hbb6fd260),
	.w3(32'h39bc8f74),
	.w4(32'hbb2cd9ea),
	.w5(32'hbc38f5db),
	.w6(32'hbaec8d52),
	.w7(32'hba377262),
	.w8(32'hbbfa9fde),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0c2df0),
	.w1(32'hbac5afd6),
	.w2(32'h3bd92bd1),
	.w3(32'hbba5e333),
	.w4(32'hbbe11ae3),
	.w5(32'h3b360be3),
	.w6(32'hbbe03f1d),
	.w7(32'hba4e24da),
	.w8(32'h3b534b74),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1b1e9f),
	.w1(32'hbb726aef),
	.w2(32'h39549e8d),
	.w3(32'h3c3c2306),
	.w4(32'hbc8e1ce9),
	.w5(32'h3b3f7d4b),
	.w6(32'h3b97b643),
	.w7(32'hbc2ff41e),
	.w8(32'hbbbc65c7),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5f59a6),
	.w1(32'h3c0f7b87),
	.w2(32'h3c889cf6),
	.w3(32'h3c323a5e),
	.w4(32'h3b72c73a),
	.w5(32'h3cb4169f),
	.w6(32'h3bbb7b9f),
	.w7(32'hbc10e339),
	.w8(32'h3cb62431),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb143f12),
	.w1(32'h3bf5fcf1),
	.w2(32'h3b8c4200),
	.w3(32'h3c5f31e1),
	.w4(32'h3b8ee0c7),
	.w5(32'h3bf36abf),
	.w6(32'h3c3d95a1),
	.w7(32'h3b7fa810),
	.w8(32'hba8204a6),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b00331b),
	.w1(32'h39b1db44),
	.w2(32'h3c382f39),
	.w3(32'h3bcdc1ac),
	.w4(32'h3bc71b3b),
	.w5(32'hbb9bb792),
	.w6(32'hbbaee9a2),
	.w7(32'h3b9709c7),
	.w8(32'h3c2eced0),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0921f6),
	.w1(32'h38ce4da5),
	.w2(32'h3c850203),
	.w3(32'hb996c9ff),
	.w4(32'h3b02dafd),
	.w5(32'h3ca72a73),
	.w6(32'h3a0d15a9),
	.w7(32'h3c1eda0e),
	.w8(32'h3c6a222b),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2e9810),
	.w1(32'h3b1b17ab),
	.w2(32'h3bb7f321),
	.w3(32'hbb55dab5),
	.w4(32'h3ba7c63b),
	.w5(32'h3c40abaa),
	.w6(32'h3b57eed3),
	.w7(32'h3b9a7113),
	.w8(32'h3be9b3a8),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b27b7eb),
	.w1(32'hbb9ccd98),
	.w2(32'hbb96f526),
	.w3(32'h3a82174d),
	.w4(32'hba24989b),
	.w5(32'hbc0596b3),
	.w6(32'h3bae8fd1),
	.w7(32'hbb1dfec9),
	.w8(32'hbbd30ea6),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb934402),
	.w1(32'hbba98304),
	.w2(32'hbb00b974),
	.w3(32'hbc0db0bb),
	.w4(32'hbb50485e),
	.w5(32'hb9bb1044),
	.w6(32'hbc036bae),
	.w7(32'hbb9e45c2),
	.w8(32'hb9d6da3f),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ada635c),
	.w1(32'h3b01248a),
	.w2(32'h3b209137),
	.w3(32'h3b886503),
	.w4(32'h3af1a913),
	.w5(32'h3b7be16f),
	.w6(32'h3b8c3d4d),
	.w7(32'h3ac12d0e),
	.w8(32'h3b3824e8),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7f483d),
	.w1(32'hbb295136),
	.w2(32'hbb4c18c0),
	.w3(32'h3a955bb1),
	.w4(32'hbb4b3afc),
	.w5(32'hba0637cc),
	.w6(32'h3b34da46),
	.w7(32'hbb1b9a5f),
	.w8(32'hbada5699),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8bc160),
	.w1(32'h3aa34783),
	.w2(32'hbb08608c),
	.w3(32'h3b905759),
	.w4(32'h3b81f5a5),
	.w5(32'hbad6d6ad),
	.w6(32'h3b3cafc6),
	.w7(32'h3b01ba73),
	.w8(32'h3ae8891d),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba6c314),
	.w1(32'h3c7fb88e),
	.w2(32'h3c8a4845),
	.w3(32'h3babf0aa),
	.w4(32'h3ccfa51f),
	.w5(32'h3cf477df),
	.w6(32'h3b2cbc05),
	.w7(32'h3c491924),
	.w8(32'h3c9625a6),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2383b7),
	.w1(32'hbaa515e0),
	.w2(32'hbb89aebb),
	.w3(32'hbb7c891a),
	.w4(32'h3bd73202),
	.w5(32'hbc181522),
	.w6(32'h3b47415f),
	.w7(32'h3aeeab9f),
	.w8(32'hbb252283),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6e587f),
	.w1(32'h3a8766fa),
	.w2(32'hba7db739),
	.w3(32'hbb7b22be),
	.w4(32'hbb778650),
	.w5(32'hbba36fac),
	.w6(32'hbb3d177f),
	.w7(32'h3bb3f615),
	.w8(32'h3b637950),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3698b71b),
	.w1(32'hbbb1ba80),
	.w2(32'h3be94e0e),
	.w3(32'hbab65745),
	.w4(32'h3b8f5709),
	.w5(32'h3c1a0f6c),
	.w6(32'hbb4d5b12),
	.w7(32'h3bf676fe),
	.w8(32'hbaaf8b63),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7fc86b),
	.w1(32'hbc1f9376),
	.w2(32'h3b0b169e),
	.w3(32'hbb2c45f1),
	.w4(32'h3909f009),
	.w5(32'h3ca69f04),
	.w6(32'hbb2075f4),
	.w7(32'h3c0b4eef),
	.w8(32'hbbad5769),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb48615a),
	.w1(32'h3b968059),
	.w2(32'h3c6b05d9),
	.w3(32'hbbd553b3),
	.w4(32'h3abff2b9),
	.w5(32'h3c3ff181),
	.w6(32'hbbd7228a),
	.w7(32'h3bf075e4),
	.w8(32'h3c283c03),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abb1d94),
	.w1(32'hbbb3ded0),
	.w2(32'hbbf601eb),
	.w3(32'h3b012bf1),
	.w4(32'hbb93e37f),
	.w5(32'hbb954248),
	.w6(32'h3bde346f),
	.w7(32'hbbc73e09),
	.w8(32'h3a5d29b8),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9b168c),
	.w1(32'hbad79627),
	.w2(32'hbc090471),
	.w3(32'h3b3b9a67),
	.w4(32'hb9153c96),
	.w5(32'h3b524f48),
	.w6(32'h3b753ed7),
	.w7(32'h3b34f8e5),
	.w8(32'h3b60b88a),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc78dc7),
	.w1(32'h3a771a5e),
	.w2(32'hbb8d516e),
	.w3(32'h3bde6ea8),
	.w4(32'hba0525e6),
	.w5(32'hb9fc33bc),
	.w6(32'h3b9a18dd),
	.w7(32'hbb37c7b7),
	.w8(32'hbbb6fe5b),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4cb0c7),
	.w1(32'hba23f99c),
	.w2(32'hbc18aa10),
	.w3(32'hbbae9ac4),
	.w4(32'h3a93008b),
	.w5(32'hbc05615c),
	.w6(32'hbb18b358),
	.w7(32'h3b491d96),
	.w8(32'hbbdc793b),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5ffd99),
	.w1(32'hbb11d8bd),
	.w2(32'hbc65f1ae),
	.w3(32'h3b109a21),
	.w4(32'hbc028c9a),
	.w5(32'hbcca2000),
	.w6(32'hba16e6c4),
	.w7(32'hbbd2d8cc),
	.w8(32'h3c2128da),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcf7311),
	.w1(32'hbbc7e30f),
	.w2(32'h3b8ef4b0),
	.w3(32'hbc11f2ff),
	.w4(32'hba0b9850),
	.w5(32'h3c197855),
	.w6(32'hbb12575c),
	.w7(32'h3b17c762),
	.w8(32'hbb56757f),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aad5cfe),
	.w1(32'h39d3b564),
	.w2(32'hbbc7a2fd),
	.w3(32'hbbb226d5),
	.w4(32'hbb832ac9),
	.w5(32'hbb403f2c),
	.w6(32'hbc3a356d),
	.w7(32'hbb7ffd24),
	.w8(32'h3b1ea505),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af3b608),
	.w1(32'h3b795176),
	.w2(32'h3c4cbe3c),
	.w3(32'h3bdd30a2),
	.w4(32'h3bca422a),
	.w5(32'h3b914ce2),
	.w6(32'h3a3b87bb),
	.w7(32'h3b43edb4),
	.w8(32'h3bbc4e1c),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3bfadf),
	.w1(32'hbba5d875),
	.w2(32'h3b3efe23),
	.w3(32'h3bd7cd4e),
	.w4(32'h3b46edb9),
	.w5(32'h3b97af8f),
	.w6(32'h3b638f39),
	.w7(32'h3b3ba30f),
	.w8(32'h3a4c5851),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39800f33),
	.w1(32'hba759349),
	.w2(32'h3c38cb79),
	.w3(32'h3b3bdd81),
	.w4(32'h39f9d5a4),
	.w5(32'h3cb0f51c),
	.w6(32'h3af54605),
	.w7(32'hba200ef2),
	.w8(32'h3a83cdb0),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb82cc9e),
	.w1(32'hbb2a45b3),
	.w2(32'h39c963c6),
	.w3(32'hba0dfbf8),
	.w4(32'hba093e96),
	.w5(32'h3c11b791),
	.w6(32'hbc2b865b),
	.w7(32'h3b9ed4bd),
	.w8(32'hbc12cf29),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b80e71c),
	.w1(32'hbc200ceb),
	.w2(32'hbbb13e13),
	.w3(32'h3bb7f5c1),
	.w4(32'hbc1de90a),
	.w5(32'hbc60f6e8),
	.w6(32'hbb24f296),
	.w7(32'hbb3c153b),
	.w8(32'hbb3b5ee9),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7e78b4),
	.w1(32'hba7f87b3),
	.w2(32'h3b0c061b),
	.w3(32'hbad7f1bd),
	.w4(32'h3a09b0d7),
	.w5(32'h3ce7af16),
	.w6(32'h3ab6c26c),
	.w7(32'h3c1e7b8b),
	.w8(32'h3b26d329),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baa0d5c),
	.w1(32'h3c1790f2),
	.w2(32'h3a2aba19),
	.w3(32'hbab02678),
	.w4(32'hbaa8f134),
	.w5(32'hbc1d8cf2),
	.w6(32'hbbd4bea6),
	.w7(32'h3b3f72bd),
	.w8(32'h3b513bb5),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc19f339),
	.w1(32'h3ba4ee3f),
	.w2(32'hbb52b539),
	.w3(32'hbb70abb0),
	.w4(32'hbc0aa814),
	.w5(32'hbc763dc1),
	.w6(32'h3a5a9690),
	.w7(32'h3aebd5d1),
	.w8(32'h3bb3d49a),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb362bf3),
	.w1(32'hbb104dc2),
	.w2(32'hbbadcc91),
	.w3(32'hbb3189e4),
	.w4(32'hbbf29696),
	.w5(32'hb9b4ae14),
	.w6(32'hbbac263a),
	.w7(32'hbb9d234e),
	.w8(32'hbae9b8e3),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b620af7),
	.w1(32'h3b6565d7),
	.w2(32'hb9871ca8),
	.w3(32'h3bed1834),
	.w4(32'h3bf42aff),
	.w5(32'h3a3fa362),
	.w6(32'h3b9862fe),
	.w7(32'hbb6acdeb),
	.w8(32'h3af1727d),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb061eb3),
	.w1(32'hba90da09),
	.w2(32'hbb884761),
	.w3(32'hbbce0b68),
	.w4(32'hbb299d0c),
	.w5(32'hbb581a1b),
	.w6(32'hbb491a8d),
	.w7(32'hbacfff58),
	.w8(32'hbb8e2b75),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae7d16e),
	.w1(32'hbb9e347f),
	.w2(32'hbbd4057a),
	.w3(32'hbb655c9d),
	.w4(32'h3b167c95),
	.w5(32'hbc19dd53),
	.w6(32'h3b218b1a),
	.w7(32'hbbfa159d),
	.w8(32'hbbb3f807),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ce46c),
	.w1(32'h3b00ac45),
	.w2(32'h3c5b855d),
	.w3(32'hbab57505),
	.w4(32'h3b8b88dc),
	.w5(32'h3c54d406),
	.w6(32'hb9c0c14d),
	.w7(32'h3c0f599b),
	.w8(32'h3c260d6f),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad3705b),
	.w1(32'h3ae87b42),
	.w2(32'h3bc91ed1),
	.w3(32'hbbde0a3c),
	.w4(32'h3bba1adf),
	.w5(32'h3b040f14),
	.w6(32'hbc216933),
	.w7(32'h3baf2efd),
	.w8(32'h3c042949),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6c0c96),
	.w1(32'hba2e0c4d),
	.w2(32'hbbcf3f42),
	.w3(32'hbb8705d2),
	.w4(32'hbc10efec),
	.w5(32'hbb9e2b90),
	.w6(32'h3958d7b4),
	.w7(32'hba38dde9),
	.w8(32'hbc40614b),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad5687b),
	.w1(32'h3aa37dcb),
	.w2(32'hbc771972),
	.w3(32'hba5ee2d5),
	.w4(32'hba846d40),
	.w5(32'hbc165b9c),
	.w6(32'hbb82cda0),
	.w7(32'hbba02238),
	.w8(32'hbc0baabb),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b818705),
	.w1(32'h3b497ebf),
	.w2(32'hbbf8581f),
	.w3(32'hbbb4018a),
	.w4(32'h3b7c02b1),
	.w5(32'hbb801c3f),
	.w6(32'hbbb8a02f),
	.w7(32'h3b792b42),
	.w8(32'hbb8b8e78),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaebf39c),
	.w1(32'h3b8e9bae),
	.w2(32'h3c3d0691),
	.w3(32'hbae3c0bd),
	.w4(32'hbb57dadb),
	.w5(32'h3b8ef40a),
	.w6(32'hbb695108),
	.w7(32'h3a0c1869),
	.w8(32'h3c2b1a3f),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b925ea7),
	.w1(32'hbb145f92),
	.w2(32'hbbac6101),
	.w3(32'hbb0ee39b),
	.w4(32'hbb30bb54),
	.w5(32'hbb2e75c2),
	.w6(32'hbb7b51ee),
	.w7(32'hbba04ec5),
	.w8(32'hbc2453b0),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8423a0),
	.w1(32'h3ba855a4),
	.w2(32'hbb023062),
	.w3(32'hbbb18ac4),
	.w4(32'hbbea8539),
	.w5(32'hbbd2d514),
	.w6(32'hbbc145cb),
	.w7(32'hbc391ce1),
	.w8(32'hbbd15491),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b283f33),
	.w1(32'h3ac0c878),
	.w2(32'hbc1f78d7),
	.w3(32'hbb26c62e),
	.w4(32'hbc39ba50),
	.w5(32'hbc0c66f3),
	.w6(32'hbb4e7ae2),
	.w7(32'h358374aa),
	.w8(32'hba13dd65),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf79f28),
	.w1(32'hbc163e24),
	.w2(32'hbc32b2fe),
	.w3(32'h3aa1f04d),
	.w4(32'hbc3c2db5),
	.w5(32'hbbb31399),
	.w6(32'h3be1742e),
	.w7(32'hbc1b1185),
	.w8(32'hbb42c909),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbb8300),
	.w1(32'h39e34f2d),
	.w2(32'hbb967f0f),
	.w3(32'hbac7cbc0),
	.w4(32'hbb6386af),
	.w5(32'h3cc95043),
	.w6(32'hb98365fc),
	.w7(32'h3afa7573),
	.w8(32'hbbeea82e),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba966e15),
	.w1(32'hbbe70694),
	.w2(32'hbb7afd3b),
	.w3(32'hbbe2ba05),
	.w4(32'h3a1f6ade),
	.w5(32'hbb90b694),
	.w6(32'hbc0cad2d),
	.w7(32'h3ba0db95),
	.w8(32'hbb8904d8),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcff58f),
	.w1(32'hbc230f6b),
	.w2(32'h3c59d91d),
	.w3(32'hbc2741dd),
	.w4(32'h3a6fcb10),
	.w5(32'h3caaeb41),
	.w6(32'hbbe0aa80),
	.w7(32'h3a0175c2),
	.w8(32'hbbd5be6b),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba7fb21),
	.w1(32'hbad70556),
	.w2(32'hb935cf35),
	.w3(32'hbc02522b),
	.w4(32'hbb818c32),
	.w5(32'h3b4c90e2),
	.w6(32'hbc805b55),
	.w7(32'hb9092c49),
	.w8(32'hb8b25902),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1a5e82),
	.w1(32'h3bf1b404),
	.w2(32'h3bf19a27),
	.w3(32'h3b5594c8),
	.w4(32'h3c98315d),
	.w5(32'h3badf84e),
	.w6(32'hbb64db21),
	.w7(32'h3bd7c8d4),
	.w8(32'hbb05b741),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd42445),
	.w1(32'hba9756d0),
	.w2(32'hbc12830a),
	.w3(32'hbc1f6f72),
	.w4(32'hbbd53510),
	.w5(32'hbc069a02),
	.w6(32'hbc4d5a98),
	.w7(32'hbbe65c8c),
	.w8(32'hbbc7fc4f),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe4e877),
	.w1(32'hba7deebc),
	.w2(32'h3afbe0c2),
	.w3(32'hbb89c65f),
	.w4(32'hba46ba5a),
	.w5(32'h3ba06c82),
	.w6(32'h3afc7868),
	.w7(32'hbbcf70b4),
	.w8(32'hbbd069ba),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9319a8),
	.w1(32'hbc4bc29b),
	.w2(32'hbc1e3751),
	.w3(32'hbb75b8ca),
	.w4(32'hbc4c6ea8),
	.w5(32'hbc958b80),
	.w6(32'hbb4afd58),
	.w7(32'hbb34558a),
	.w8(32'hbc58b342),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3e4b11),
	.w1(32'hbbf4c4f4),
	.w2(32'hbbaf3ab7),
	.w3(32'h3b2b210c),
	.w4(32'h397c8bd1),
	.w5(32'hbb01f264),
	.w6(32'hbbcaecf5),
	.w7(32'hbb6ede89),
	.w8(32'hbbd90804),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf6b9a1),
	.w1(32'h3a9750a7),
	.w2(32'hbaf47395),
	.w3(32'hbb86b92f),
	.w4(32'hbb9cc1c6),
	.w5(32'h3b976767),
	.w6(32'hb9e1d0a7),
	.w7(32'hbaa9b76a),
	.w8(32'h3c13bc79),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4088d4),
	.w1(32'h3bccab5c),
	.w2(32'hbb521e55),
	.w3(32'h39c21cab),
	.w4(32'h3b3c2cf7),
	.w5(32'hbb0fc466),
	.w6(32'hba722c8e),
	.w7(32'hbb831348),
	.w8(32'h3bdedd9a),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad9817d),
	.w1(32'h3b91dded),
	.w2(32'hbadac683),
	.w3(32'h3b849763),
	.w4(32'h3aacdb65),
	.w5(32'h3cd23374),
	.w6(32'h3c029ed2),
	.w7(32'hbb3e351b),
	.w8(32'hbb8d3782),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc32685c),
	.w1(32'hbc310350),
	.w2(32'h3bfa6d87),
	.w3(32'hbc88c19c),
	.w4(32'hbbbb370f),
	.w5(32'h3c1fb55d),
	.w6(32'hbb9d62c3),
	.w7(32'hba04b9ca),
	.w8(32'hb992a79a),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd9abdb),
	.w1(32'hbba578b2),
	.w2(32'hbbbe6c12),
	.w3(32'hbb1309d0),
	.w4(32'hbbf5eb66),
	.w5(32'hbb5e55e7),
	.w6(32'hbb2e8355),
	.w7(32'hb9aaeb6e),
	.w8(32'hb9cf86c4),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf71d64),
	.w1(32'h3ae7b6ae),
	.w2(32'hbabd7593),
	.w3(32'hbb303b84),
	.w4(32'h3ac947f0),
	.w5(32'hbc612d82),
	.w6(32'h3b02f78d),
	.w7(32'hbafe8735),
	.w8(32'hbb3012b3),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8bc991),
	.w1(32'h3b537c6d),
	.w2(32'h3aed9218),
	.w3(32'h3b3b094e),
	.w4(32'h3ba3b470),
	.w5(32'hbb6a8904),
	.w6(32'hb9c7a036),
	.w7(32'hbb35fd60),
	.w8(32'hbb0a21a0),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf91ee4),
	.w1(32'hbc19dbe5),
	.w2(32'hbbee21e7),
	.w3(32'hbc6f8005),
	.w4(32'hbc1a955c),
	.w5(32'hbca3fae9),
	.w6(32'hbb399f62),
	.w7(32'hbbc65106),
	.w8(32'hbb434a60),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbbb964),
	.w1(32'hbb3fb925),
	.w2(32'h3c5ce909),
	.w3(32'hbc58aae0),
	.w4(32'h3a469e4c),
	.w5(32'h3d00f354),
	.w6(32'hbb122a20),
	.w7(32'h3bb469dc),
	.w8(32'h3b9f0e6b),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe0ed1f),
	.w1(32'hbacacab7),
	.w2(32'h3ba53557),
	.w3(32'hbc06cfa2),
	.w4(32'hbb415ae7),
	.w5(32'h3b93fec0),
	.w6(32'hbb89f1cd),
	.w7(32'hba296ee3),
	.w8(32'h3b0556a9),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb67d30a2),
	.w1(32'hbb026552),
	.w2(32'hbab23613),
	.w3(32'h3bc2d5ac),
	.w4(32'hbbb38833),
	.w5(32'h3ada8d32),
	.w6(32'hbb39df41),
	.w7(32'hbbe37ecb),
	.w8(32'hbbdc3b2d),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2c8299),
	.w1(32'h3c0a0b8b),
	.w2(32'hbb14f565),
	.w3(32'hbb0e71ee),
	.w4(32'h3ba1115f),
	.w5(32'h3b94599b),
	.w6(32'hbb218f4f),
	.w7(32'h3b5de7f5),
	.w8(32'hbba097d6),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba31dbbb),
	.w1(32'hbc2546af),
	.w2(32'hbc4ef1c8),
	.w3(32'h3ae291ee),
	.w4(32'hbc2086e3),
	.w5(32'hbc1f083b),
	.w6(32'h3b350d89),
	.w7(32'hbc0e06cc),
	.w8(32'h3b74dc45),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b78f7e4),
	.w1(32'hbae0477d),
	.w2(32'hbb76e192),
	.w3(32'h3c682fb5),
	.w4(32'hbb9ee9aa),
	.w5(32'hbc21c933),
	.w6(32'h3c2bb7e2),
	.w7(32'hbb28a08b),
	.w8(32'hba3e2ee2),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a126a8b),
	.w1(32'hbc293652),
	.w2(32'h3c271781),
	.w3(32'hb9c34226),
	.w4(32'h3a707787),
	.w5(32'h3d041e1e),
	.w6(32'hbab62b03),
	.w7(32'hbb661181),
	.w8(32'hbc1c91d7),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4c34ed),
	.w1(32'hbbf5f3de),
	.w2(32'hbc0ec8d9),
	.w3(32'hbbfcf1b7),
	.w4(32'hbbf1c8d7),
	.w5(32'hbbb5fe60),
	.w6(32'hbb9d654e),
	.w7(32'hbb2608dc),
	.w8(32'hbbaab14e),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb997ecad),
	.w1(32'hbc5238cc),
	.w2(32'hbbacd685),
	.w3(32'hbb5b6ffe),
	.w4(32'hbbb3603b),
	.w5(32'h3c13c6ad),
	.w6(32'h3b1a6244),
	.w7(32'h3b8752e4),
	.w8(32'hbbdc28f7),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule