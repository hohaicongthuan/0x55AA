module layer_10_featuremap_59(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398a3bba),
	.w1(32'h3ab44598),
	.w2(32'hba3b0c9f),
	.w3(32'h381076ba),
	.w4(32'h3a83d0fa),
	.w5(32'h3a4143e5),
	.w6(32'hbb388f27),
	.w7(32'hbab9bad1),
	.w8(32'h3ae87522),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb492b8d),
	.w1(32'h3b8544e7),
	.w2(32'h3c4ab9b0),
	.w3(32'h3ada00cf),
	.w4(32'h3b3dd217),
	.w5(32'h3b30dec0),
	.w6(32'h3b21d23d),
	.w7(32'h3b524b2c),
	.w8(32'h3b2f5e17),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2fe63d),
	.w1(32'hbb2d69b7),
	.w2(32'hb8ca167a),
	.w3(32'hbb408e9a),
	.w4(32'hbb549f95),
	.w5(32'h3a7aa61d),
	.w6(32'hbb0c696e),
	.w7(32'hbae0de01),
	.w8(32'hba39be07),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafc2576),
	.w1(32'hba9f3284),
	.w2(32'h3a97e8c6),
	.w3(32'h3937b861),
	.w4(32'h3a190108),
	.w5(32'h3b1929f0),
	.w6(32'hbb1b4cc7),
	.w7(32'hba9822ac),
	.w8(32'hbab750f8),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b118370),
	.w1(32'h3a339ffe),
	.w2(32'h3b6ec856),
	.w3(32'h3b03bb70),
	.w4(32'hbac2312b),
	.w5(32'h3b34e96b),
	.w6(32'hbade0416),
	.w7(32'hbb874f25),
	.w8(32'h3b080755),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98bd419),
	.w1(32'h3a98d3c6),
	.w2(32'h3ab0fbfd),
	.w3(32'hbab46289),
	.w4(32'h39f38291),
	.w5(32'h3a7e8c23),
	.w6(32'hbb04794d),
	.w7(32'h3a45e8d0),
	.w8(32'h3a1d5bc2),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6c5d47),
	.w1(32'h3b8c381a),
	.w2(32'hbc97c771),
	.w3(32'h3b6cc5ea),
	.w4(32'h3bbcc44f),
	.w5(32'hb9a5d16a),
	.w6(32'h3b068a5c),
	.w7(32'h3b9ce7fc),
	.w8(32'h3bac1586),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8be1e3),
	.w1(32'h3b56b40a),
	.w2(32'h3cb933a3),
	.w3(32'h3d571b94),
	.w4(32'h3ca75d88),
	.w5(32'h3bf120a6),
	.w6(32'h3cc088a2),
	.w7(32'hbae75345),
	.w8(32'hbc685d69),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb55e85e),
	.w1(32'hbaf69425),
	.w2(32'h3b036f73),
	.w3(32'hbb279175),
	.w4(32'hbb031989),
	.w5(32'h38bac44c),
	.w6(32'hbb5c0b99),
	.w7(32'hbb2c1098),
	.w8(32'h39b88abf),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8a0950),
	.w1(32'hbbfeb726),
	.w2(32'hbc857dd9),
	.w3(32'hbc12c3b7),
	.w4(32'hbc369ced),
	.w5(32'hbbbfd876),
	.w6(32'hba8a80eb),
	.w7(32'hbb9e5353),
	.w8(32'h3bff7072),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5bb88a),
	.w1(32'h39e89375),
	.w2(32'hba10c0a3),
	.w3(32'h3a1cb048),
	.w4(32'h39c66dd8),
	.w5(32'h3abc60db),
	.w6(32'h3a244ce2),
	.w7(32'h399899bd),
	.w8(32'h3aaba1e5),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1b1b59),
	.w1(32'h3b97595d),
	.w2(32'hbcc31b68),
	.w3(32'hbb81f66e),
	.w4(32'h391f75f0),
	.w5(32'hbc387e14),
	.w6(32'h3a50a443),
	.w7(32'h3bf4ca61),
	.w8(32'h3ca6c76c),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb238a92),
	.w1(32'hbbf66386),
	.w2(32'hbc65380b),
	.w3(32'hba8dd227),
	.w4(32'hbb442aba),
	.w5(32'hbb707f8f),
	.w6(32'hbba197ca),
	.w7(32'hbb634c6c),
	.w8(32'h39522146),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b78abbd),
	.w1(32'hbb97f705),
	.w2(32'h39a4a314),
	.w3(32'h3b8c217e),
	.w4(32'h3b228e53),
	.w5(32'h3b4fe357),
	.w6(32'h3bb34771),
	.w7(32'hbb36949c),
	.w8(32'h3996f9e5),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9b5033),
	.w1(32'h3c2853b6),
	.w2(32'h3ba7cc7d),
	.w3(32'hb9c66713),
	.w4(32'hba8fb46a),
	.w5(32'hbba207a3),
	.w6(32'h3b165eff),
	.w7(32'h3b98429c),
	.w8(32'h3ad2082a),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca00bd4),
	.w1(32'hbc9df22e),
	.w2(32'hbc9954dd),
	.w3(32'hbc120af8),
	.w4(32'hbc3265b3),
	.w5(32'hbb2541dd),
	.w6(32'h3c328eb8),
	.w7(32'h3bb04187),
	.w8(32'h3bb9bab4),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ecbacd),
	.w1(32'hba317bac),
	.w2(32'h3a6594c6),
	.w3(32'hba233849),
	.w4(32'hba04918e),
	.w5(32'hba08e6df),
	.w6(32'hb93129e3),
	.w7(32'hb9eaf7a2),
	.w8(32'hbb48483f),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac24f3d),
	.w1(32'hbc1987bc),
	.w2(32'hbcca2ca2),
	.w3(32'h3cac433f),
	.w4(32'h3bb067a6),
	.w5(32'h3c1c751a),
	.w6(32'hbbacfe1d),
	.w7(32'hba8c20a0),
	.w8(32'h3b5c4857),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba83efde),
	.w1(32'hbba2093b),
	.w2(32'hbc94835c),
	.w3(32'h3bc1351d),
	.w4(32'h395a02b9),
	.w5(32'hbaf451b8),
	.w6(32'hbb9cd3d0),
	.w7(32'hbb3f8642),
	.w8(32'hbb8eebfe),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaecc393),
	.w1(32'hbb00935f),
	.w2(32'h398cebb4),
	.w3(32'h39f7001e),
	.w4(32'hba66bb8c),
	.w5(32'hb8d5d3d0),
	.w6(32'hbab1b046),
	.w7(32'hbab3b3a1),
	.w8(32'hb9f6746f),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba166137),
	.w1(32'h3a1fe6ea),
	.w2(32'h3ac5d356),
	.w3(32'hba744e2f),
	.w4(32'h3a980bda),
	.w5(32'h3b4674e2),
	.w6(32'hba6659fa),
	.w7(32'h3a294fe2),
	.w8(32'h37729454),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae3b126),
	.w1(32'h3b4dd28a),
	.w2(32'h3b1389e8),
	.w3(32'hba0187a7),
	.w4(32'hba6bc487),
	.w5(32'hba584272),
	.w6(32'hbae1ed27),
	.w7(32'hbaf303b2),
	.w8(32'hbad7d1dc),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b880110),
	.w1(32'hbc70e6b8),
	.w2(32'hbd1906a9),
	.w3(32'h3cebdacb),
	.w4(32'h3aa372cf),
	.w5(32'hbb141651),
	.w6(32'h3d0b1315),
	.w7(32'hbc0789a7),
	.w8(32'h3c20c32c),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9864189),
	.w1(32'h3a25a9bb),
	.w2(32'hbac70bfa),
	.w3(32'hba63bd6e),
	.w4(32'hbb1c20f5),
	.w5(32'hbbbb84e7),
	.w6(32'hb732a31d),
	.w7(32'h3a18c8ed),
	.w8(32'h3b3a168a),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc90be9a),
	.w1(32'h3c6b4cb7),
	.w2(32'h3cba1b6d),
	.w3(32'hbc95cfad),
	.w4(32'hbb6a2877),
	.w5(32'hbba5460a),
	.w6(32'hbc8f454c),
	.w7(32'hbbc28123),
	.w8(32'hbbef5770),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b48821e),
	.w1(32'h3b1e7ec2),
	.w2(32'hbb27504b),
	.w3(32'h3abad38b),
	.w4(32'h3a04440d),
	.w5(32'hba57bfd0),
	.w6(32'hba778379),
	.w7(32'hbaf9f10c),
	.w8(32'hbaeeb2dc),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa0cde6),
	.w1(32'hb99d87de),
	.w2(32'hb80873e7),
	.w3(32'h39233bfe),
	.w4(32'h3ac9abb2),
	.w5(32'hb9d286d5),
	.w6(32'hbad10775),
	.w7(32'hba76df8b),
	.w8(32'hba484d2c),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd6f1412),
	.w1(32'h3c59958b),
	.w2(32'h3b095896),
	.w3(32'hbd5b1e78),
	.w4(32'hbbd6317f),
	.w5(32'hbc74d5b5),
	.w6(32'hbd064b4e),
	.w7(32'h3c613a2a),
	.w8(32'h3c827fc0),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc51b9d),
	.w1(32'hbba7bba5),
	.w2(32'h3b0bd165),
	.w3(32'hbc090ac2),
	.w4(32'hbb7847b2),
	.w5(32'hb9fe8f59),
	.w6(32'hbb8db7ea),
	.w7(32'hbb1df714),
	.w8(32'hbc504b4f),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1f58fd),
	.w1(32'hba99c77f),
	.w2(32'h3b1cf725),
	.w3(32'hbd5bd660),
	.w4(32'hbcf6bf52),
	.w5(32'hbc92b204),
	.w6(32'hbd150f5d),
	.w7(32'hbafb7305),
	.w8(32'hbc2dd825),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb994d37),
	.w1(32'hbacec8b3),
	.w2(32'h3bc1ce8f),
	.w3(32'hbb0a172a),
	.w4(32'hba5a67e1),
	.w5(32'h3c7e9fcb),
	.w6(32'hbb27efa8),
	.w7(32'hbb658229),
	.w8(32'hbc13d6b4),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a175d97),
	.w1(32'hbb7eb924),
	.w2(32'h3c61e39b),
	.w3(32'hbc2cf032),
	.w4(32'hbbe34135),
	.w5(32'h3b3992be),
	.w6(32'hbc474ebb),
	.w7(32'h399f192d),
	.w8(32'hbc8d5cd4),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1b3f09),
	.w1(32'hbc1cf1d2),
	.w2(32'hba29d6b0),
	.w3(32'hbb3a2f16),
	.w4(32'hbc12f740),
	.w5(32'h3bdc1e89),
	.w6(32'h3b7cd354),
	.w7(32'h3c45ff4c),
	.w8(32'h3ba72ff8),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb14c700),
	.w1(32'h3bd5a2ef),
	.w2(32'h3c15f4fc),
	.w3(32'hba8c49ba),
	.w4(32'h3b39d74b),
	.w5(32'hbbc3a895),
	.w6(32'hbb96e759),
	.w7(32'hbb8ae857),
	.w8(32'hbbeb7d1b),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf4fe04),
	.w1(32'h3a888226),
	.w2(32'hbb8d3e19),
	.w3(32'h3baa7c2e),
	.w4(32'h3c09eb9b),
	.w5(32'h3ad408a2),
	.w6(32'h3c157f8a),
	.w7(32'hbb5fa652),
	.w8(32'h3afe4675),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba41328),
	.w1(32'h3b2959ca),
	.w2(32'hbc0b8c15),
	.w3(32'h3c2310db),
	.w4(32'h3bcee853),
	.w5(32'h3c21dfc5),
	.w6(32'hbb35e303),
	.w7(32'hbc15656c),
	.w8(32'hb94aaaaa),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d45fb6f),
	.w1(32'h3cafb051),
	.w2(32'hbc0431b9),
	.w3(32'h3cc20caa),
	.w4(32'hbc2958d0),
	.w5(32'hbd0c6df4),
	.w6(32'h3c877d47),
	.w7(32'hbca6128b),
	.w8(32'h3c0a7eaa),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc89f2b7),
	.w1(32'h3cced185),
	.w2(32'h3cf77e49),
	.w3(32'hbd122b46),
	.w4(32'hbc6d258b),
	.w5(32'hbcdd7b89),
	.w6(32'hbd0d80c4),
	.w7(32'hbc371722),
	.w8(32'hbbc35383),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1d9bf9),
	.w1(32'h3c6f5442),
	.w2(32'h3cdbc79c),
	.w3(32'hbd4cf328),
	.w4(32'h3b9cc68f),
	.w5(32'hbb89bb5e),
	.w6(32'hbc80dd10),
	.w7(32'h3c7b1db4),
	.w8(32'h3c6794d6),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b29f945),
	.w1(32'hbac031c8),
	.w2(32'h3b8fa622),
	.w3(32'h3b304822),
	.w4(32'hbc2fb00c),
	.w5(32'hbb8dedfa),
	.w6(32'hbb03f0e6),
	.w7(32'hbacc7371),
	.w8(32'hbb38ba66),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb42fdd2),
	.w1(32'h3ba3ac2a),
	.w2(32'h3b28f55c),
	.w3(32'hbb927b96),
	.w4(32'h39efd96a),
	.w5(32'hbb00b889),
	.w6(32'hbbaeb575),
	.w7(32'hbb1de009),
	.w8(32'hbb0ca61f),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba97b138),
	.w1(32'hbb61ed48),
	.w2(32'h3c6655a5),
	.w3(32'h3ac726aa),
	.w4(32'h3b815f6b),
	.w5(32'hbc55e4d8),
	.w6(32'h3c0a55e4),
	.w7(32'h3ae22170),
	.w8(32'hbca06e72),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0626b6),
	.w1(32'hbc244ce0),
	.w2(32'h3afed475),
	.w3(32'hbcb7f284),
	.w4(32'hbb32adcc),
	.w5(32'hbafffa05),
	.w6(32'h3bc7dcc8),
	.w7(32'h3c835f87),
	.w8(32'h3a67d5ab),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd91650),
	.w1(32'hbc8bdda4),
	.w2(32'hbc3df8e6),
	.w3(32'hbc9d396a),
	.w4(32'hbc66d8c1),
	.w5(32'h3cb3a79a),
	.w6(32'hbc584dd8),
	.w7(32'h3afb6b2f),
	.w8(32'h3c43109e),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba02b2d8),
	.w1(32'h3b2fde9e),
	.w2(32'hbba7b019),
	.w3(32'hbcf0e9bc),
	.w4(32'hbd1d6da1),
	.w5(32'hbca90c3d),
	.w6(32'hbcc41f03),
	.w7(32'hbc50dac3),
	.w8(32'hbb219f7e),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b22a8d5),
	.w1(32'h3c8ad55c),
	.w2(32'h38e839c4),
	.w3(32'h3b991bf6),
	.w4(32'h3c30f70e),
	.w5(32'hbbddbc2e),
	.w6(32'h3cfdaac6),
	.w7(32'h3c8fc145),
	.w8(32'h3c21fb4a),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc843929),
	.w1(32'h3bb1ecaf),
	.w2(32'hbb264176),
	.w3(32'h3c1f9abc),
	.w4(32'h3bacc3f8),
	.w5(32'hbbc660c5),
	.w6(32'h3c2e81fc),
	.w7(32'hbb9b3675),
	.w8(32'h3ba96bb1),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c92c8ae),
	.w1(32'hbc9bd4a2),
	.w2(32'hbd1ba0e1),
	.w3(32'h3cfc5f44),
	.w4(32'h3bc17ef8),
	.w5(32'hbba52121),
	.w6(32'h3c17babf),
	.w7(32'hbc65552e),
	.w8(32'hbafde463),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3911b6d2),
	.w1(32'hbb107e48),
	.w2(32'h3c289c51),
	.w3(32'hbaf3ba87),
	.w4(32'hbb0cdd5e),
	.w5(32'hba9d8297),
	.w6(32'hba56355e),
	.w7(32'hbb042129),
	.w8(32'hbc390fd7),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc145740),
	.w1(32'h3c201174),
	.w2(32'h3a384b0e),
	.w3(32'hbc4f193f),
	.w4(32'h3c8b4144),
	.w5(32'hbc41d0e2),
	.w6(32'h3a9ea355),
	.w7(32'h3ba4c229),
	.w8(32'h391cf8d2),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae4e3ab),
	.w1(32'h3b39e7d9),
	.w2(32'h3ae9def4),
	.w3(32'hbb8f6853),
	.w4(32'hbb94b030),
	.w5(32'hbb457a95),
	.w6(32'hbc176f52),
	.w7(32'h3b472ff2),
	.w8(32'hbbb8006e),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf8f599),
	.w1(32'hbc40a106),
	.w2(32'hbb707bff),
	.w3(32'hbcbc93fd),
	.w4(32'hbb1d3037),
	.w5(32'h3b105105),
	.w6(32'hbc443fd0),
	.w7(32'h3bce3410),
	.w8(32'hbaa16a03),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a015691),
	.w1(32'hbb8ab41d),
	.w2(32'h3b7ae732),
	.w3(32'h3c188cd5),
	.w4(32'h3aaa312a),
	.w5(32'h390c44bb),
	.w6(32'hbb1e294b),
	.w7(32'h3bac1f89),
	.w8(32'hba0c641c),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5df423),
	.w1(32'hbcadb382),
	.w2(32'hbcf703aa),
	.w3(32'h3bf1a2e8),
	.w4(32'hbb6cc5bf),
	.w5(32'h3c027c39),
	.w6(32'h3af29bd2),
	.w7(32'hbbbb80b5),
	.w8(32'h3c75366a),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba6c67c),
	.w1(32'hb9850e36),
	.w2(32'h3c15b316),
	.w3(32'h3a48036e),
	.w4(32'hbc7383b4),
	.w5(32'h3cfe7d2d),
	.w6(32'hbca28290),
	.w7(32'hbc6412d7),
	.w8(32'h3abcfcfc),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9312ec),
	.w1(32'h3bba5ee0),
	.w2(32'hbc01dfed),
	.w3(32'h3cc10a07),
	.w4(32'hbc0ea663),
	.w5(32'hbb7c8a85),
	.w6(32'hbcab516b),
	.w7(32'hbb4d8200),
	.w8(32'h3c9fd051),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb029b57),
	.w1(32'h3a696198),
	.w2(32'h3b5e9ea4),
	.w3(32'h3c52cd72),
	.w4(32'hbc15a312),
	.w5(32'h3b705d16),
	.w6(32'h3b3b46cf),
	.w7(32'hbc47831e),
	.w8(32'h3b8fdaf4),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1d8d9e),
	.w1(32'h3b457007),
	.w2(32'hbb284b39),
	.w3(32'hbb638f73),
	.w4(32'hb92ab9e7),
	.w5(32'hbb7b5a11),
	.w6(32'hbb9c03f4),
	.w7(32'h3b1d2d2e),
	.w8(32'hbc34b32f),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4a859d),
	.w1(32'h3b85da9d),
	.w2(32'h3b2ebe64),
	.w3(32'hba956cd9),
	.w4(32'h39b9f984),
	.w5(32'h3b0f6966),
	.w6(32'hbbd243fd),
	.w7(32'hbb890cac),
	.w8(32'h3ad7eecd),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8bdfa5),
	.w1(32'hbb6abcc8),
	.w2(32'hbb034baf),
	.w3(32'h38605eb0),
	.w4(32'h3b0feafd),
	.w5(32'hbbc1e288),
	.w6(32'h3a1d7d4d),
	.w7(32'hba990181),
	.w8(32'h3afe3b87),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc28065c),
	.w1(32'hbb1e86b3),
	.w2(32'hbc96503c),
	.w3(32'hbb882ba5),
	.w4(32'h3bfa7ff2),
	.w5(32'hbc45faa7),
	.w6(32'hbaaf283b),
	.w7(32'h3ba9917b),
	.w8(32'h3b572589),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd36d11b),
	.w1(32'hbc2768d6),
	.w2(32'hbcb90026),
	.w3(32'h3b0ab8a6),
	.w4(32'h3c1f3a8e),
	.w5(32'hbc7b4996),
	.w6(32'h3c040280),
	.w7(32'h3c0ba477),
	.w8(32'h3bf3cca3),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc689fe6),
	.w1(32'h380006fe),
	.w2(32'hba77e06c),
	.w3(32'hba8d1ce6),
	.w4(32'h3c83122f),
	.w5(32'hbb67aa41),
	.w6(32'h3c8a7539),
	.w7(32'h3c5012b1),
	.w8(32'h3ad7aa9b),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb605a49),
	.w1(32'hbaa961d3),
	.w2(32'hbb30e560),
	.w3(32'hbad98719),
	.w4(32'hbb676b56),
	.w5(32'h3cceb53e),
	.w6(32'h3a450d93),
	.w7(32'h3a954ecc),
	.w8(32'h3bd819f4),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfa0fc5),
	.w1(32'hbb15d774),
	.w2(32'h3b342593),
	.w3(32'h3c2e448b),
	.w4(32'h3b36b6fc),
	.w5(32'h3b4e7d2a),
	.w6(32'hbbd1f61b),
	.w7(32'hbbf36dd3),
	.w8(32'hbb1697e2),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a314d69),
	.w1(32'hbb34ac9a),
	.w2(32'h3b690439),
	.w3(32'hba023456),
	.w4(32'hbbb4c692),
	.w5(32'h3b5c206d),
	.w6(32'hbb4c5fea),
	.w7(32'hbb744ca1),
	.w8(32'h3bdf04b5),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd03eca),
	.w1(32'hbd27ad87),
	.w2(32'hbd40c5c0),
	.w3(32'hbc9d6394),
	.w4(32'hbcdaa578),
	.w5(32'hbb8a368e),
	.w6(32'h3cf0e537),
	.w7(32'h3cb974a1),
	.w8(32'h3d33c691),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb004529),
	.w1(32'hbc41492b),
	.w2(32'h3c0129bb),
	.w3(32'h3c911147),
	.w4(32'h3a83f1c1),
	.w5(32'h3cbfad18),
	.w6(32'hbd08a1d1),
	.w7(32'hbcc7b0c3),
	.w8(32'hbb6533a6),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7f604b),
	.w1(32'hbb620b5b),
	.w2(32'hbc54df94),
	.w3(32'h3c00771b),
	.w4(32'h3bc40d16),
	.w5(32'h3c3273d9),
	.w6(32'hbb70be3b),
	.w7(32'h3b1d0f76),
	.w8(32'hbbbe76ed),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce79c2c),
	.w1(32'h3c9721fe),
	.w2(32'h3d095999),
	.w3(32'hbd10d6d8),
	.w4(32'hbc799202),
	.w5(32'hbc34d683),
	.w6(32'hbd15a57f),
	.w7(32'hbc288dc3),
	.w8(32'hbc09445c),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a38e8d8),
	.w1(32'hbb89ebf9),
	.w2(32'h3b66fe18),
	.w3(32'hbbab538b),
	.w4(32'hbc24d334),
	.w5(32'h3a85da7d),
	.w6(32'hbb2fb32d),
	.w7(32'hbc0e2701),
	.w8(32'h3bb0e3c1),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5e116d),
	.w1(32'h39d6c79a),
	.w2(32'hbbf27f1d),
	.w3(32'h3b0bd7c8),
	.w4(32'h3ba03724),
	.w5(32'h3c4163f0),
	.w6(32'h3aba658d),
	.w7(32'h3b8b2980),
	.w8(32'h3ba365df),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ad999f),
	.w1(32'h3c1ad6dc),
	.w2(32'h3c1dc78c),
	.w3(32'h3c4b4b65),
	.w4(32'hbc2e95c6),
	.w5(32'hbc0c1465),
	.w6(32'hbc1eb266),
	.w7(32'hbd24b4f2),
	.w8(32'hbc25242c),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc196ec7),
	.w1(32'hbc986030),
	.w2(32'hbc00b759),
	.w3(32'hbcf3b12c),
	.w4(32'h3b0f99d3),
	.w5(32'hbb1e5a74),
	.w6(32'hbc15e47c),
	.w7(32'h3d0bf5da),
	.w8(32'hbb79e6be),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2bca63),
	.w1(32'hba9456ca),
	.w2(32'h3b09abcf),
	.w3(32'hbb01f334),
	.w4(32'hbacea9fe),
	.w5(32'hbb8efa53),
	.w6(32'h3a844334),
	.w7(32'hbae91cdd),
	.w8(32'hb9f4d60a),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4f7e0c),
	.w1(32'hbb45d37d),
	.w2(32'hbcec35d6),
	.w3(32'h3a8c49bb),
	.w4(32'h3b1bc9a8),
	.w5(32'h3b13151e),
	.w6(32'h3b1388f5),
	.w7(32'hba3a1118),
	.w8(32'h3c7fc672),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c346a76),
	.w1(32'hbbec2496),
	.w2(32'hbcc00c24),
	.w3(32'h3d0c6b8a),
	.w4(32'h3bf4c08e),
	.w5(32'h3c58da4c),
	.w6(32'h3c2e818c),
	.w7(32'hbc8d110e),
	.w8(32'h3bb4fd74),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc37b06a),
	.w1(32'h3b75bced),
	.w2(32'hbb9f5d39),
	.w3(32'hbc5128d7),
	.w4(32'hbc985c8c),
	.w5(32'hbc89c491),
	.w6(32'hbc75ecd4),
	.w7(32'hbc536d27),
	.w8(32'h3b490ee2),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0139c4),
	.w1(32'hba3dee9d),
	.w2(32'hbbee2734),
	.w3(32'h3baf9146),
	.w4(32'hbad32da7),
	.w5(32'h3ba51949),
	.w6(32'h3c391e09),
	.w7(32'hbba0f3d0),
	.w8(32'h3b468170),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9b0461),
	.w1(32'hbc08311e),
	.w2(32'hbca9504e),
	.w3(32'hbac654d4),
	.w4(32'hbc5053aa),
	.w5(32'hbc01f91b),
	.w6(32'h3c122988),
	.w7(32'h3c22c325),
	.w8(32'h3ca43f23),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc24bbba),
	.w1(32'h3a845c4e),
	.w2(32'hb9ae16d9),
	.w3(32'hbc91c930),
	.w4(32'hbbdce716),
	.w5(32'hbb772153),
	.w6(32'hbc120176),
	.w7(32'hba088b30),
	.w8(32'h3a4cb51c),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5e1748),
	.w1(32'hbabc68d6),
	.w2(32'hbcac902b),
	.w3(32'h3b1b6f20),
	.w4(32'h394fec76),
	.w5(32'hbc7a57d1),
	.w6(32'hbae29828),
	.w7(32'hbb0af909),
	.w8(32'h3bf779bf),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc89bd33),
	.w1(32'hba9bdcfa),
	.w2(32'hbb5724ad),
	.w3(32'h3ccccf69),
	.w4(32'h3ca7563b),
	.w5(32'hbc353d7a),
	.w6(32'h3ce8ce87),
	.w7(32'hbc181239),
	.w8(32'hbc0e0186),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbac12e2),
	.w1(32'hbb0e24b1),
	.w2(32'hbc84129f),
	.w3(32'h3b8a77c3),
	.w4(32'hbb35320d),
	.w5(32'hbb4a075c),
	.w6(32'h3b86f3fd),
	.w7(32'hb94b0628),
	.w8(32'h3cbf1232),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb364731),
	.w1(32'h3c710d8e),
	.w2(32'h3c0aa0bf),
	.w3(32'h3caff78a),
	.w4(32'h3c68ae05),
	.w5(32'h3c340d3c),
	.w6(32'h3ca43878),
	.w7(32'hbc81479e),
	.w8(32'h3ab12ae6),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39dea46f),
	.w1(32'hbc095ba4),
	.w2(32'h3aa239ab),
	.w3(32'hbc157e57),
	.w4(32'hbc5f325d),
	.w5(32'hba6e115c),
	.w6(32'hbcc54b96),
	.w7(32'hbb09c8fd),
	.w8(32'hbb76e679),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe0b605),
	.w1(32'h3c4efc1b),
	.w2(32'h3c605199),
	.w3(32'hbc7e13f4),
	.w4(32'hbac3c34b),
	.w5(32'hbbbbc556),
	.w6(32'hbc1ab8b1),
	.w7(32'h3b703d12),
	.w8(32'h3b769a9f),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5c708c),
	.w1(32'hbaf1806d),
	.w2(32'h3a8e5b97),
	.w3(32'hbb41006a),
	.w4(32'hba7e724d),
	.w5(32'hbc1ab785),
	.w6(32'h3ad902d8),
	.w7(32'h3ad83329),
	.w8(32'hbc0ce62b),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd1a2c5),
	.w1(32'h38e812be),
	.w2(32'h3c260a68),
	.w3(32'hb9f60d83),
	.w4(32'h3b0f8196),
	.w5(32'h3c3498d4),
	.w6(32'hbc075950),
	.w7(32'h3c16cf83),
	.w8(32'hbb37589f),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8994f0),
	.w1(32'hbc43afb3),
	.w2(32'hbc3dc87b),
	.w3(32'h3c8b94ed),
	.w4(32'h3ad3c1da),
	.w5(32'hbb010743),
	.w6(32'h3a86ca45),
	.w7(32'hbc1709a3),
	.w8(32'hbbdf1716),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4532cb),
	.w1(32'h3bb79d10),
	.w2(32'h3bbc6615),
	.w3(32'hbcbed5ad),
	.w4(32'hbb78b31d),
	.w5(32'hbbef4721),
	.w6(32'hbc30cc70),
	.w7(32'h3c146bef),
	.w8(32'h3b6176e4),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc45503),
	.w1(32'hbcb3bbc2),
	.w2(32'hbd64d61f),
	.w3(32'hbb859df8),
	.w4(32'hbc8a31d7),
	.w5(32'hbd081340),
	.w6(32'h3d1d9e45),
	.w7(32'h3ba43d11),
	.w8(32'h3c49371a),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f5a301),
	.w1(32'h3c7e8aea),
	.w2(32'h3c170110),
	.w3(32'hbc9c6397),
	.w4(32'hbb634f83),
	.w5(32'hbbbf95c5),
	.w6(32'hbc8dbdd3),
	.w7(32'hbb8ed4ad),
	.w8(32'hb95edc74),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc82ab21),
	.w1(32'hbc5e726a),
	.w2(32'hbcb55b2f),
	.w3(32'h3bc01810),
	.w4(32'hba7c0ceb),
	.w5(32'h3b6bacb9),
	.w6(32'h3c2fb59b),
	.w7(32'h3b6520a2),
	.w8(32'h3c25ec6c),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4ad6d7),
	.w1(32'hbc38ee6c),
	.w2(32'hbb68f037),
	.w3(32'hbc1192b1),
	.w4(32'hbc25f53c),
	.w5(32'hbc511f66),
	.w6(32'h3c33c1a4),
	.w7(32'h3c58d059),
	.w8(32'hba450211),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb26ecf),
	.w1(32'h3b38e501),
	.w2(32'h3c10690c),
	.w3(32'hbd135059),
	.w4(32'h3a26a046),
	.w5(32'hbcba3f09),
	.w6(32'hbc209933),
	.w7(32'h3c300596),
	.w8(32'hbb39671f),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb852ec5),
	.w1(32'hbb0f8d89),
	.w2(32'hbcbf9ed5),
	.w3(32'hbc74cbd3),
	.w4(32'hbc418806),
	.w5(32'hbd032459),
	.w6(32'hbbde5871),
	.w7(32'hbc48cb84),
	.w8(32'h3c15f57a),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8b1303),
	.w1(32'h3baf8f77),
	.w2(32'hbc9015fd),
	.w3(32'h3cfa6695),
	.w4(32'h3cffb775),
	.w5(32'h3be3576c),
	.w6(32'h3d0f7596),
	.w7(32'h3c64f63c),
	.w8(32'h3bc18422),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be0e0e3),
	.w1(32'hbc8bb208),
	.w2(32'hbd1f3f08),
	.w3(32'hbcd1ef1f),
	.w4(32'hbca8039b),
	.w5(32'hbd00b21a),
	.w6(32'h3b9f0626),
	.w7(32'h3c25caee),
	.w8(32'h3cbfd794),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c016caa),
	.w1(32'h3c681bf8),
	.w2(32'h3c993039),
	.w3(32'h3c1abe72),
	.w4(32'hbbe708e8),
	.w5(32'hbbf3e656),
	.w6(32'h3c9a061b),
	.w7(32'hbd1dec83),
	.w8(32'hbcdf905d),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb118b9),
	.w1(32'h3c38ec27),
	.w2(32'h3d301193),
	.w3(32'hbd2f1803),
	.w4(32'hbc0dc620),
	.w5(32'h3cc280fb),
	.w6(32'hbc9c27b8),
	.w7(32'h3c584da2),
	.w8(32'h39bf050a),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb71abf4),
	.w1(32'h3b98d83f),
	.w2(32'h3c29816a),
	.w3(32'hbc9394b3),
	.w4(32'hbc8d242f),
	.w5(32'hbc59fff3),
	.w6(32'hbd107531),
	.w7(32'hb9d043f0),
	.w8(32'hbc657e2b),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5af944),
	.w1(32'hbcb8e377),
	.w2(32'hbd1669fe),
	.w3(32'h3b40fb41),
	.w4(32'hbc9affad),
	.w5(32'hbcbbdf45),
	.w6(32'h3d05afff),
	.w7(32'hbc102f67),
	.w8(32'h3c3e4ef8),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9b4d9a),
	.w1(32'h3b4829c5),
	.w2(32'h3ba3a256),
	.w3(32'hbc2ca67c),
	.w4(32'h3b2292fa),
	.w5(32'h3b7d403a),
	.w6(32'hbb98b00d),
	.w7(32'h3b530fd7),
	.w8(32'hbb310d3a),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d09df8e),
	.w1(32'h3caa97db),
	.w2(32'hbbd22cb0),
	.w3(32'h3c8ab901),
	.w4(32'h3c5fff97),
	.w5(32'hbce19400),
	.w6(32'h3c45651e),
	.w7(32'hbd05b8eb),
	.w8(32'hbc92cc97),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf3f1f9),
	.w1(32'h3afc78a1),
	.w2(32'hbb4f8da2),
	.w3(32'hbc5aee2e),
	.w4(32'h3b705159),
	.w5(32'hbbd0e44c),
	.w6(32'hbb5833ff),
	.w7(32'h3b1fb9f9),
	.w8(32'hbb4df121),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb58b7f1),
	.w1(32'hbb6a7404),
	.w2(32'hbb553910),
	.w3(32'hbbd5997d),
	.w4(32'hbb8bd47a),
	.w5(32'hbb3e7c0e),
	.w6(32'hbc345cf7),
	.w7(32'hbb8264bd),
	.w8(32'hbb19ea2f),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6c2960),
	.w1(32'hbb0a5715),
	.w2(32'hbc9f2164),
	.w3(32'hbad07954),
	.w4(32'hbbb85138),
	.w5(32'h3b71f36f),
	.w6(32'h3b6f2981),
	.w7(32'hb98ed20a),
	.w8(32'h3ca16dcf),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8f74f8),
	.w1(32'hbb443663),
	.w2(32'h3768a121),
	.w3(32'h3c1f1438),
	.w4(32'hbb4a3167),
	.w5(32'hbb5d36ff),
	.w6(32'hbbdea12f),
	.w7(32'hbcdab5a5),
	.w8(32'hbc73e138),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbfbf02),
	.w1(32'h3b0ac576),
	.w2(32'h3aefcdad),
	.w3(32'hbcdfa017),
	.w4(32'hbc1adcb1),
	.w5(32'hbcdb6446),
	.w6(32'hbcb72cd8),
	.w7(32'h3c7c7fe0),
	.w8(32'hbbb2642c),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcab11c2),
	.w1(32'h3c0211af),
	.w2(32'h3c0860fb),
	.w3(32'hbc9e0688),
	.w4(32'h3c18aff5),
	.w5(32'hbc11b15a),
	.w6(32'h3c141359),
	.w7(32'h3d03a721),
	.w8(32'h3b8b28ee),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba478c64),
	.w1(32'h3c1ee413),
	.w2(32'h3b5fb852),
	.w3(32'h3afd7e5d),
	.w4(32'h3b67d374),
	.w5(32'hbc242b48),
	.w6(32'hbbead358),
	.w7(32'hbb903e41),
	.w8(32'h3b9a26cf),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc935fd5),
	.w1(32'h3c4178d5),
	.w2(32'h3cb90ed0),
	.w3(32'h3c57331b),
	.w4(32'h3d187bf9),
	.w5(32'hbc048f3c),
	.w6(32'h3c213d1c),
	.w7(32'hbb543545),
	.w8(32'hbd03c0f1),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3852d4),
	.w1(32'hbcdc2a77),
	.w2(32'hbc6b8991),
	.w3(32'hbbe5cacb),
	.w4(32'hbc1e8dfa),
	.w5(32'hb810844e),
	.w6(32'h3cf018fc),
	.w7(32'h3cd8a51c),
	.w8(32'h3c75e95d),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb24ad4),
	.w1(32'h3beb1af1),
	.w2(32'h3baf16e8),
	.w3(32'hbbfb3170),
	.w4(32'hbc173766),
	.w5(32'h3b719cd7),
	.w6(32'hbc74f9ee),
	.w7(32'hbbe265d8),
	.w8(32'h3b49f8e7),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2a55ba),
	.w1(32'h3aa9e82b),
	.w2(32'h3bd013f5),
	.w3(32'h3b2e84cb),
	.w4(32'h3aef148d),
	.w5(32'h3b6de15e),
	.w6(32'hbae0591f),
	.w7(32'hbbec0630),
	.w8(32'hb9362047),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adcf510),
	.w1(32'h3a80a379),
	.w2(32'h3af0d02d),
	.w3(32'h3b60ac56),
	.w4(32'hbb005f39),
	.w5(32'h3b70a7e4),
	.w6(32'h3a0eded4),
	.w7(32'hbafa6cd6),
	.w8(32'h399315bb),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb30a895),
	.w1(32'hbb9541df),
	.w2(32'h3a05be60),
	.w3(32'h3b06035a),
	.w4(32'h3b0d6c11),
	.w5(32'h3c63cf01),
	.w6(32'h3a147dc8),
	.w7(32'hbaf124aa),
	.w8(32'hbb70fed6),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aefde1f),
	.w1(32'h3ab37a1f),
	.w2(32'h3c86f58d),
	.w3(32'hbbd2df51),
	.w4(32'hbc081fd8),
	.w5(32'h3c99ff56),
	.w6(32'hbc8b174a),
	.w7(32'hbab6e94c),
	.w8(32'hbbb9d5be),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc052c0a),
	.w1(32'hbbf0121b),
	.w2(32'h3b4bcc62),
	.w3(32'hbc6a2f54),
	.w4(32'hbc1eb00e),
	.w5(32'hbcb3193a),
	.w6(32'hbcb0d389),
	.w7(32'h3babcd8d),
	.w8(32'hbc47640a),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc860f51),
	.w1(32'hbbcec8bd),
	.w2(32'hbb898931),
	.w3(32'hbcc11138),
	.w4(32'h3babbde5),
	.w5(32'hbb72a87f),
	.w6(32'hba2535ca),
	.w7(32'h3cab3af9),
	.w8(32'hbb0bfdd4),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b37c61e),
	.w1(32'hbbca260d),
	.w2(32'hbc430ffc),
	.w3(32'h3b618ae9),
	.w4(32'hbb378971),
	.w5(32'hbbc28521),
	.w6(32'h3b963fa3),
	.w7(32'h3a0a7101),
	.w8(32'h3b1cf424),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8afb5f),
	.w1(32'h3c238afc),
	.w2(32'h3c6a8112),
	.w3(32'hbc48cef6),
	.w4(32'hbb2b1e0a),
	.w5(32'hbbc67b15),
	.w6(32'hbc757b00),
	.w7(32'hbb936726),
	.w8(32'hba652f4d),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb929fe0),
	.w1(32'hbbe18f46),
	.w2(32'h3a3fac9c),
	.w3(32'hbbd1e3dd),
	.w4(32'h3c0b9cd4),
	.w5(32'hba14e7f4),
	.w6(32'h3a64d59d),
	.w7(32'h3bd1d2d7),
	.w8(32'h3ac1db88),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb367b57),
	.w1(32'hbabbaed5),
	.w2(32'hba8691c4),
	.w3(32'hba28685e),
	.w4(32'h3b5418b7),
	.w5(32'h3928417f),
	.w6(32'h3b2b1ef3),
	.w7(32'h3b411968),
	.w8(32'hbbffc932),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b03bb2a),
	.w1(32'hbb92cb2c),
	.w2(32'hbb5b074e),
	.w3(32'h3a2e4e80),
	.w4(32'hbbdec17f),
	.w5(32'h3aef4080),
	.w6(32'hbc1d822a),
	.w7(32'hbbf79402),
	.w8(32'hbc346345),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad83cb5),
	.w1(32'h3ab334f4),
	.w2(32'h3b70a08c),
	.w3(32'h3b884612),
	.w4(32'hbc47ab09),
	.w5(32'h3c6375fa),
	.w6(32'hbcc28a7b),
	.w7(32'hbccd3deb),
	.w8(32'hbbff796e),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c587b08),
	.w1(32'hbb872e9f),
	.w2(32'h3c2eff88),
	.w3(32'h3caedf24),
	.w4(32'h3be8a8c9),
	.w5(32'h3c02de53),
	.w6(32'hbd25bb7e),
	.w7(32'hbd4b6ec5),
	.w8(32'h3b03c6b0),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb33e74c),
	.w1(32'hbc06d3d6),
	.w2(32'hbce06ed0),
	.w3(32'h3bc4a3eb),
	.w4(32'hbc0eb606),
	.w5(32'hbc7de708),
	.w6(32'h3c7afc14),
	.w7(32'h3ac2f13e),
	.w8(32'h3c5814d9),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb55ed68),
	.w1(32'h3bb8b586),
	.w2(32'hbb8215d4),
	.w3(32'hbaea577e),
	.w4(32'h3c1f9fba),
	.w5(32'hbb6489d4),
	.w6(32'h3cbc130e),
	.w7(32'h3c173330),
	.w8(32'hbb570649),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc374490),
	.w1(32'hbc4c62d5),
	.w2(32'h3c5c66da),
	.w3(32'hbb661df2),
	.w4(32'h3c259ed6),
	.w5(32'hbc03fe4f),
	.w6(32'h3b30789f),
	.w7(32'h3b7089c1),
	.w8(32'hbcb2bbd8),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc26dab9),
	.w1(32'hbc17724c),
	.w2(32'hbbd8fc7d),
	.w3(32'hbcb51672),
	.w4(32'h3a9bd6ab),
	.w5(32'hbc1822fc),
	.w6(32'h399c3678),
	.w7(32'h3cb6994b),
	.w8(32'h3b13627d),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeba5e8),
	.w1(32'hb7c1ffd2),
	.w2(32'h3c661d98),
	.w3(32'hbb51f75d),
	.w4(32'h3ad45768),
	.w5(32'h3cd1e339),
	.w6(32'h3b3e2fdf),
	.w7(32'h3ae429f1),
	.w8(32'h39da2729),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb22d9e3),
	.w1(32'hbbf5a3fa),
	.w2(32'hbbbb51bd),
	.w3(32'hbc68a1ad),
	.w4(32'hbcc25be6),
	.w5(32'hbc0c2fc6),
	.w6(32'hbcc6d58a),
	.w7(32'hbaee2530),
	.w8(32'h3b861366),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0e9a45),
	.w1(32'hbc4f110f),
	.w2(32'hbcc8de7e),
	.w3(32'h3c180bde),
	.w4(32'hbb043dd7),
	.w5(32'h3bbe091f),
	.w6(32'h3b407551),
	.w7(32'h3a58fcef),
	.w8(32'h3bbcc18b),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af6297b),
	.w1(32'h3b67f77f),
	.w2(32'h3c1c1e14),
	.w3(32'hbbaa7480),
	.w4(32'hb94cb50a),
	.w5(32'hbb8926ef),
	.w6(32'hbbdab7b5),
	.w7(32'hbb90f191),
	.w8(32'hbae8219c),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1cfa55),
	.w1(32'hbc6e99d8),
	.w2(32'hbb8e0fa2),
	.w3(32'h3ba1a487),
	.w4(32'hbc1a710a),
	.w5(32'h3baaca58),
	.w6(32'h3bbd3b75),
	.w7(32'hbbdd5f10),
	.w8(32'h3be80c23),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5f180f),
	.w1(32'hbbe6e780),
	.w2(32'hbcd22770),
	.w3(32'h3c55bdb2),
	.w4(32'h3900d873),
	.w5(32'hbb7cb1ae),
	.w6(32'h3b2499fe),
	.w7(32'hbb7bc5d4),
	.w8(32'h3b67dfe8),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbee4824),
	.w1(32'h3bd0661e),
	.w2(32'h3d0bdf65),
	.w3(32'hbb7b24ad),
	.w4(32'h3b0972ad),
	.w5(32'hbae885e4),
	.w6(32'hbba657da),
	.w7(32'hbbf57fdb),
	.w8(32'hbcb1538f),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf3c413),
	.w1(32'hbc4e0995),
	.w2(32'hbc86d252),
	.w3(32'hbce8da1a),
	.w4(32'hbc1bdc92),
	.w5(32'hbbe95bea),
	.w6(32'h3a0582fa),
	.w7(32'h3ca45077),
	.w8(32'h3bd023b9),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb817858),
	.w1(32'hb90d2399),
	.w2(32'hbb423aa6),
	.w3(32'hbb29dd12),
	.w4(32'hbad8dbc7),
	.w5(32'hba893cbc),
	.w6(32'hbb005cc5),
	.w7(32'hbac4edd8),
	.w8(32'h3a0687a3),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce9b1ab),
	.w1(32'h3c513d32),
	.w2(32'h3c856027),
	.w3(32'hbd04c550),
	.w4(32'h3b334a6d),
	.w5(32'hbc1c7d3a),
	.w6(32'hbc60906b),
	.w7(32'h3bf0defe),
	.w8(32'h3b366179),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beeecd0),
	.w1(32'h3c2e35f0),
	.w2(32'h3bdfc732),
	.w3(32'hbae91e54),
	.w4(32'h3c2bc926),
	.w5(32'h3c1b9eeb),
	.w6(32'h3c082c4f),
	.w7(32'hbbb82b29),
	.w8(32'h3ba263ac),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2bce3a),
	.w1(32'hbbab6ce2),
	.w2(32'hbae61cde),
	.w3(32'hbb2abb93),
	.w4(32'hba9ca8bc),
	.w5(32'hba42f038),
	.w6(32'hbb536ba1),
	.w7(32'hbaaf5b42),
	.w8(32'hb91ca927),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb917e40b),
	.w1(32'h3b42d707),
	.w2(32'hbac430df),
	.w3(32'h3a6a0e70),
	.w4(32'h3b748467),
	.w5(32'hbb4e2a2e),
	.w6(32'h3aaeeaf6),
	.w7(32'h3a978751),
	.w8(32'hba20db54),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc205bec),
	.w1(32'hbb60c27b),
	.w2(32'hbad1e99f),
	.w3(32'hbc5c39d0),
	.w4(32'hbbb87658),
	.w5(32'hbc0016cc),
	.w6(32'h3c05aec1),
	.w7(32'h3c0d5de8),
	.w8(32'h3c28af5d),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a630ed4),
	.w1(32'h3c657675),
	.w2(32'hba702b02),
	.w3(32'hba842e54),
	.w4(32'h3a4751c9),
	.w5(32'hbc9e74dd),
	.w6(32'h3b3f69e2),
	.w7(32'h3bfb82da),
	.w8(32'h3a107bb2),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc588f1d),
	.w1(32'hbc1fd99b),
	.w2(32'hbbd48653),
	.w3(32'hbb058db7),
	.w4(32'h3baba548),
	.w5(32'h3afd95c9),
	.w6(32'h3bf54380),
	.w7(32'h3c077baa),
	.w8(32'h3b192b8b),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa20189),
	.w1(32'h3b991200),
	.w2(32'hbca17255),
	.w3(32'hbb54c133),
	.w4(32'h3ad2941f),
	.w5(32'hbce4a10d),
	.w6(32'hbb41d732),
	.w7(32'h3b91acd3),
	.w8(32'h3c2b747a),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca665e8),
	.w1(32'hba1c3ef2),
	.w2(32'hbc783b6d),
	.w3(32'h3b977de1),
	.w4(32'h3cb902f6),
	.w5(32'hbc02ba65),
	.w6(32'h3d0aa194),
	.w7(32'h3c914a6a),
	.w8(32'h3b893555),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba50c8d),
	.w1(32'hbb9628d7),
	.w2(32'hbaedfb1b),
	.w3(32'hbb714285),
	.w4(32'h3abc76d3),
	.w5(32'hba4015f9),
	.w6(32'hba65a266),
	.w7(32'h3b9a112a),
	.w8(32'h399c3f10),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c15ad94),
	.w1(32'hbca222d9),
	.w2(32'hbd094f47),
	.w3(32'h3c27648d),
	.w4(32'hbc5d9b54),
	.w5(32'hbc4d9704),
	.w6(32'h3ca1eb83),
	.w7(32'hb9e3a8d8),
	.w8(32'h3b64f25c),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcdbff19),
	.w1(32'h3c1e7085),
	.w2(32'h3bd8fb9d),
	.w3(32'hbd3f155b),
	.w4(32'hbcaf2e83),
	.w5(32'hbd0b92a4),
	.w6(32'hbd37f4af),
	.w7(32'hbbfddd7e),
	.w8(32'h3b09752b),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3fb4e1),
	.w1(32'h3c65bdc2),
	.w2(32'h389b3135),
	.w3(32'h3921b7f4),
	.w4(32'h3d0771a6),
	.w5(32'h3c61db31),
	.w6(32'h3cfaed8e),
	.w7(32'h3cbb7a68),
	.w8(32'h3c0ee22d),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9de5058),
	.w1(32'h3b2715ff),
	.w2(32'hbb00a094),
	.w3(32'h3b414636),
	.w4(32'hbaa9db29),
	.w5(32'hbb1af9cf),
	.w6(32'hba87908b),
	.w7(32'h3bafd06f),
	.w8(32'hba888c85),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfc51b1),
	.w1(32'h3ad1b70b),
	.w2(32'h3c8686fd),
	.w3(32'hbc23a6ec),
	.w4(32'hbb824c9b),
	.w5(32'h3bc4dd71),
	.w6(32'hbc135c4a),
	.w7(32'hba9b8cdc),
	.w8(32'h3a4153a3),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0c7d24),
	.w1(32'h3cc8ea1c),
	.w2(32'h3a897baf),
	.w3(32'hbc15869a),
	.w4(32'h3a84a6f1),
	.w5(32'hbc1f006a),
	.w6(32'hbbcf9b7c),
	.w7(32'h3c4db8f8),
	.w8(32'h3bce01a6),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc359a05),
	.w1(32'h3c25ef2e),
	.w2(32'h3bc6c3e2),
	.w3(32'hbbe78d15),
	.w4(32'hbb93066a),
	.w5(32'hbb5dfed1),
	.w6(32'h3c3c7a97),
	.w7(32'h3be49413),
	.w8(32'hbadf2a54),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbc909e),
	.w1(32'hbb3400d7),
	.w2(32'hbc1d794a),
	.w3(32'h3bebd74b),
	.w4(32'hbb3b2284),
	.w5(32'hbba9370a),
	.w6(32'h3bc51e74),
	.w7(32'hbb3e4254),
	.w8(32'h3b152e97),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad49402),
	.w1(32'hbae77e66),
	.w2(32'hba41e943),
	.w3(32'h3c9f41ae),
	.w4(32'h3c654b74),
	.w5(32'hba4d8649),
	.w6(32'h3cb8496c),
	.w7(32'h3c5ac9bf),
	.w8(32'h3a8cdb50),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c62a82c),
	.w1(32'hbb515c38),
	.w2(32'hbbb42727),
	.w3(32'h3c44b7c9),
	.w4(32'h3c383af8),
	.w5(32'h3c13f8b9),
	.w6(32'h3c98914f),
	.w7(32'h3c0727fe),
	.w8(32'h3bc34993),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c20948c),
	.w1(32'h3ba60518),
	.w2(32'hbbeea96d),
	.w3(32'h3b4ed1d1),
	.w4(32'h3ababdcf),
	.w5(32'hbb70dcb6),
	.w6(32'h3a92869b),
	.w7(32'hba4e42b4),
	.w8(32'h3985869e),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc42ef7c),
	.w1(32'h3b1ffd6e),
	.w2(32'h3c3243ff),
	.w3(32'hbb53a932),
	.w4(32'h3c5b8812),
	.w5(32'h3af1edaa),
	.w6(32'hbcd0400c),
	.w7(32'hbc97961d),
	.w8(32'hba2a1942),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b21be0b),
	.w1(32'h3b3d4fcd),
	.w2(32'h3a625fd7),
	.w3(32'hbb9b8ce7),
	.w4(32'h3acf9e74),
	.w5(32'h3bd33efc),
	.w6(32'hbb75e7de),
	.w7(32'hb92de626),
	.w8(32'hbaf2d933),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b99b799),
	.w1(32'hbb15d241),
	.w2(32'h3bf507bf),
	.w3(32'h3cbb4230),
	.w4(32'h3cb8afd9),
	.w5(32'h3b642568),
	.w6(32'hbc12aaf4),
	.w7(32'hbbacffd0),
	.w8(32'hba95662e),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3935bb),
	.w1(32'h3c123fa7),
	.w2(32'hbb5c5932),
	.w3(32'hbacac1f9),
	.w4(32'hbbf2948b),
	.w5(32'h3b014526),
	.w6(32'hbb5040a2),
	.w7(32'hbc18ae2a),
	.w8(32'hbc3b6df9),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c512c9f),
	.w1(32'h3c01837a),
	.w2(32'h388e8deb),
	.w3(32'h3b1a21b5),
	.w4(32'hbac57a94),
	.w5(32'hbbe71a8a),
	.w6(32'hbc3e0ea0),
	.w7(32'hbc07f8ce),
	.w8(32'h3ba51471),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf9e7c4),
	.w1(32'h3c764ede),
	.w2(32'hba8cc7a2),
	.w3(32'hbcbc84c6),
	.w4(32'hbba7f3be),
	.w5(32'hbc082617),
	.w6(32'hbb8e0ccd),
	.w7(32'h3ba0377c),
	.w8(32'hbb9aa66e),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1f11e6),
	.w1(32'hbc3f3ea2),
	.w2(32'h3bcffe32),
	.w3(32'h3b7abf6b),
	.w4(32'h3b2fe2e3),
	.w5(32'h3c57ef5e),
	.w6(32'hbc575065),
	.w7(32'hbc9252d4),
	.w8(32'hbc197e2b),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca9e6c4),
	.w1(32'h3c9cb55d),
	.w2(32'h3b498589),
	.w3(32'h3ce090f2),
	.w4(32'h3ceb894d),
	.w5(32'h3a174f76),
	.w6(32'hbc024da7),
	.w7(32'h3bf34320),
	.w8(32'h3b67164d),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4dfdf2),
	.w1(32'hbbc29821),
	.w2(32'h3c206669),
	.w3(32'hbb2b2cef),
	.w4(32'h3b8c5b53),
	.w5(32'hbb645388),
	.w6(32'hbbacc858),
	.w7(32'hbc31aa51),
	.w8(32'hbb488a3e),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4342fa),
	.w1(32'hba09f865),
	.w2(32'hbbeac777),
	.w3(32'hbc930a7e),
	.w4(32'hbba26608),
	.w5(32'hbcaac8e1),
	.w6(32'hbc135c00),
	.w7(32'h3bbc9610),
	.w8(32'hbb976788),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce9d3fa),
	.w1(32'hbc98d463),
	.w2(32'hbc845328),
	.w3(32'hbce92ca8),
	.w4(32'hbca9223a),
	.w5(32'hbc31330a),
	.w6(32'hbca0ea30),
	.w7(32'h3bb6994e),
	.w8(32'h3b812118),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6161e0),
	.w1(32'h3ab55e5f),
	.w2(32'hbc90b170),
	.w3(32'hbb1de9e1),
	.w4(32'hbb15e56a),
	.w5(32'hbb2841ca),
	.w6(32'h3c9ab93c),
	.w7(32'h3bb1af3c),
	.w8(32'h3b8331c8),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc85888e),
	.w1(32'hbc350f0b),
	.w2(32'hbc7f4d1a),
	.w3(32'hbc02f4f2),
	.w4(32'hbbb32402),
	.w5(32'h3a33bae0),
	.w6(32'hbb253f0b),
	.w7(32'hbb2739c0),
	.w8(32'h3bb4514a),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0fc82b),
	.w1(32'hbc5142fb),
	.w2(32'h3bc70850),
	.w3(32'hbb8103f9),
	.w4(32'h39c204bb),
	.w5(32'hb7e2c082),
	.w6(32'hbbe9bd51),
	.w7(32'h3b1015b6),
	.w8(32'h3b81e0c8),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2732a3),
	.w1(32'hbbb445be),
	.w2(32'hbc99c979),
	.w3(32'hbbc2541b),
	.w4(32'hbb2d3e26),
	.w5(32'h3c27b5c8),
	.w6(32'h3b8685b3),
	.w7(32'h3c1eeb41),
	.w8(32'h3ca13c0a),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f0914d),
	.w1(32'hbb5f82bb),
	.w2(32'h3b0009b8),
	.w3(32'h3b49a2d4),
	.w4(32'hbb85f2e1),
	.w5(32'h3b5a9671),
	.w6(32'h3c462ca4),
	.w7(32'hbb41186c),
	.w8(32'hbc19e76c),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d0c51d7),
	.w1(32'h3cbe723d),
	.w2(32'hbb5bef1a),
	.w3(32'h3ccf4fe9),
	.w4(32'h3ca0c264),
	.w5(32'hbc29e1d9),
	.w6(32'h3bc55c8b),
	.w7(32'h3ad4bf70),
	.w8(32'hbc887f6d),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc0112f),
	.w1(32'h3c666735),
	.w2(32'h3c1e978b),
	.w3(32'h3bf84d10),
	.w4(32'h3be2deb5),
	.w5(32'h3c03a834),
	.w6(32'hbc0cf513),
	.w7(32'hbc829244),
	.w8(32'hbc40ecb5),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c11e182),
	.w1(32'h3c2b58d4),
	.w2(32'hbcfe9659),
	.w3(32'h3cd11c2e),
	.w4(32'h3c083c70),
	.w5(32'hbc4cac21),
	.w6(32'h3c44bd0f),
	.w7(32'h3b94b705),
	.w8(32'hbbbc705c),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd310d0),
	.w1(32'hbb09fce6),
	.w2(32'h3af21c52),
	.w3(32'h3c17f824),
	.w4(32'h3bce1a77),
	.w5(32'h3b72ff72),
	.w6(32'hbba147d3),
	.w7(32'hbb73d1de),
	.w8(32'hb9d28980),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf3674f),
	.w1(32'h3c5249cc),
	.w2(32'h3a87ac56),
	.w3(32'h3c99aa98),
	.w4(32'h3c58e775),
	.w5(32'hbbc949e6),
	.w6(32'h3ad9942e),
	.w7(32'hba8d6fdb),
	.w8(32'hbb01dc2f),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe7b09b),
	.w1(32'hbb364b9a),
	.w2(32'hbb9a56fc),
	.w3(32'hbc61d1ff),
	.w4(32'h363fded0),
	.w5(32'hbc856e3b),
	.w6(32'h392077ce),
	.w7(32'hbb59e386),
	.w8(32'hbbb679be),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6b3a10),
	.w1(32'hbb60d1f4),
	.w2(32'hbca24f2d),
	.w3(32'hbc40531e),
	.w4(32'hbc465cf3),
	.w5(32'hbbc0a11e),
	.w6(32'h3880f599),
	.w7(32'hbb9eca87),
	.w8(32'hbbe7a964),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c61de80),
	.w1(32'h3c20f037),
	.w2(32'h3a5df5a6),
	.w3(32'hbb264e08),
	.w4(32'h3b21b457),
	.w5(32'hbc7573f8),
	.w6(32'hbb1c9a30),
	.w7(32'hbbe47ac8),
	.w8(32'h3b80ae77),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4e20de),
	.w1(32'hbc0f1bbb),
	.w2(32'hbc0bb016),
	.w3(32'hbb2a90c8),
	.w4(32'hbc0171c6),
	.w5(32'hbbcc07e1),
	.w6(32'h3b94426d),
	.w7(32'hbb535400),
	.w8(32'hbc1971f7),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc76aa0b),
	.w1(32'hbca9630f),
	.w2(32'hbcc8300a),
	.w3(32'h3c08ef5d),
	.w4(32'h3aff8ba3),
	.w5(32'h3c95582d),
	.w6(32'hbccb0952),
	.w7(32'hbc7c9f59),
	.w8(32'h3c5254ea),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd526536),
	.w1(32'h393388b0),
	.w2(32'hbbd323ee),
	.w3(32'hbd32b076),
	.w4(32'hbc9f0287),
	.w5(32'hbca5e555),
	.w6(32'hbc5f6a7f),
	.w7(32'h3c8735e5),
	.w8(32'h3c979740),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaf5b3e),
	.w1(32'h3b180712),
	.w2(32'hbc123a5c),
	.w3(32'hba081c7a),
	.w4(32'hba4858c4),
	.w5(32'hba62424e),
	.w6(32'h3c9fadb8),
	.w7(32'h3bb01c60),
	.w8(32'h3c66ea31),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc1c7c3),
	.w1(32'h3c03c557),
	.w2(32'h3b4405d4),
	.w3(32'h3c155afc),
	.w4(32'h3c73a220),
	.w5(32'h3b56e226),
	.w6(32'h3c94d339),
	.w7(32'h3c79056a),
	.w8(32'hbc735f50),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c28012a),
	.w1(32'h3b61c65e),
	.w2(32'h3b873775),
	.w3(32'h3c28b4cf),
	.w4(32'hba9ee763),
	.w5(32'h38f81c42),
	.w6(32'hbc68898f),
	.w7(32'hbcbb74dc),
	.w8(32'h3ba5b73b),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe8ee60),
	.w1(32'hbc1d6a54),
	.w2(32'hbbf320f9),
	.w3(32'hbc06747b),
	.w4(32'hbc26ddeb),
	.w5(32'hbbdd3946),
	.w6(32'h3a9895e2),
	.w7(32'h3b8cc4be),
	.w8(32'hba60c181),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae3b692),
	.w1(32'h3b33d9fd),
	.w2(32'h3a453244),
	.w3(32'hbac3d37d),
	.w4(32'h3b43b5f1),
	.w5(32'h3adac2e0),
	.w6(32'h395c279c),
	.w7(32'h39d16acc),
	.w8(32'hb9319adc),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c131ab3),
	.w1(32'h3bbb0c4a),
	.w2(32'h3c424276),
	.w3(32'h3b1bc178),
	.w4(32'h3a746ad8),
	.w5(32'h3c7513e1),
	.w6(32'hbb112c09),
	.w7(32'hbb504d61),
	.w8(32'hbb8bbdaa),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8174b8),
	.w1(32'h3bed4b01),
	.w2(32'h3ca33455),
	.w3(32'h3bd157d3),
	.w4(32'h3b016831),
	.w5(32'hbc0febd4),
	.w6(32'hb9e88617),
	.w7(32'hba40702a),
	.w8(32'hbbc4d586),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7c9afa),
	.w1(32'h3ca4d0a7),
	.w2(32'hbc0abdb9),
	.w3(32'h3bf55667),
	.w4(32'h3c6a45eb),
	.w5(32'hbc1aafdf),
	.w6(32'hbb8e35cf),
	.w7(32'h3a0d6a86),
	.w8(32'hbc0c942b),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1422f4),
	.w1(32'hbc918ffd),
	.w2(32'hbbe51571),
	.w3(32'hbc20ad87),
	.w4(32'hbc3e3714),
	.w5(32'h3b98628d),
	.w6(32'hbc6e003b),
	.w7(32'hbc729850),
	.w8(32'h3be0c128),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab850ca),
	.w1(32'h3aba1834),
	.w2(32'hbb997663),
	.w3(32'h372910b4),
	.w4(32'hbb14cfd9),
	.w5(32'hbbd73209),
	.w6(32'h3a40b363),
	.w7(32'hbba907d0),
	.w8(32'h3a335b9d),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc076b88),
	.w1(32'hba94b0b2),
	.w2(32'hbb7f9422),
	.w3(32'hba788c46),
	.w4(32'hbb1e6d67),
	.w5(32'h3b996500),
	.w6(32'h3bbe729b),
	.w7(32'h3b659a3e),
	.w8(32'h3c28bcb5),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc543b58),
	.w1(32'hbc8e3819),
	.w2(32'hbc81708a),
	.w3(32'hbbc5e989),
	.w4(32'h3acb4b3b),
	.w5(32'hbca321ca),
	.w6(32'h3c17a0c6),
	.w7(32'h3950eed0),
	.w8(32'hbbcc1734),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd577e6),
	.w1(32'h3c3ebebf),
	.w2(32'h3bd88ad2),
	.w3(32'h3b9142d6),
	.w4(32'h3c23e4e3),
	.w5(32'hba1ae2e4),
	.w6(32'hbbeea474),
	.w7(32'hbbba9fef),
	.w8(32'h3b935a46),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a586891),
	.w1(32'h3b14cf60),
	.w2(32'hbbe61770),
	.w3(32'hbb8d2910),
	.w4(32'h3ad1e882),
	.w5(32'hbba0b41c),
	.w6(32'hbb4f0881),
	.w7(32'h3b3440af),
	.w8(32'hbb8ea879),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc05137a),
	.w1(32'h3c1b857d),
	.w2(32'h3c6decee),
	.w3(32'hbc9a1673),
	.w4(32'hbc466605),
	.w5(32'hbc82d919),
	.w6(32'hbc237c2f),
	.w7(32'hbb57d694),
	.w8(32'hbb9d18e8),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc070647),
	.w1(32'h3b2a96e0),
	.w2(32'hbb3935b3),
	.w3(32'hbc0fd28f),
	.w4(32'hbb28ae12),
	.w5(32'hbbc0763d),
	.w6(32'hbbb9d67d),
	.w7(32'hbb50b297),
	.w8(32'hba4864a3),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb92e802),
	.w1(32'h3b4bdb8f),
	.w2(32'h3a940df2),
	.w3(32'h3c8d0413),
	.w4(32'h3c854333),
	.w5(32'h3a8ea79c),
	.w6(32'hbbf78699),
	.w7(32'hbbbeae81),
	.w8(32'h3b100b09),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc89c5eb),
	.w1(32'hba8a77de),
	.w2(32'h3bd33f21),
	.w3(32'hbca399b5),
	.w4(32'hbc393be6),
	.w5(32'hbc04a5dc),
	.w6(32'hba662adb),
	.w7(32'h3c3674ea),
	.w8(32'h3a8e6f50),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc25dc6f),
	.w1(32'hbbe62423),
	.w2(32'hbbe90b8e),
	.w3(32'hbc2686d7),
	.w4(32'hbc09747c),
	.w5(32'h3aba4deb),
	.w6(32'hbb300ab2),
	.w7(32'hbb811f2a),
	.w8(32'hbaf69c63),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc049a02),
	.w1(32'hbbcc7e4a),
	.w2(32'hb8f458ce),
	.w3(32'hbb5c9441),
	.w4(32'h37955886),
	.w5(32'hbb0531e2),
	.w6(32'hbc6c8edd),
	.w7(32'hbc28ceaa),
	.w8(32'h3a7682f3),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b739f28),
	.w1(32'h3b6ad03d),
	.w2(32'h3b1bc51a),
	.w3(32'hbab76abb),
	.w4(32'hbb45c01e),
	.w5(32'h3c32ddbd),
	.w6(32'hba6ce02c),
	.w7(32'hbaacd87d),
	.w8(32'h3bde0279),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ad1a4b),
	.w1(32'hbc4c06cf),
	.w2(32'h3a9d4838),
	.w3(32'h3b0085c6),
	.w4(32'hbcbf9051),
	.w5(32'h3b4c237b),
	.w6(32'hbbfa511a),
	.w7(32'hbc23fc54),
	.w8(32'h3bca700c),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bb047e),
	.w1(32'hbb234f9a),
	.w2(32'h3c87461e),
	.w3(32'h3b268bb2),
	.w4(32'hbb61dfe2),
	.w5(32'h3c5586e2),
	.w6(32'hbc24eeba),
	.w7(32'hbc896fcf),
	.w8(32'h3c2838f2),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7d1842),
	.w1(32'h39851584),
	.w2(32'hbbe97759),
	.w3(32'h3c8c37b9),
	.w4(32'h3c0d642f),
	.w5(32'h3c63b095),
	.w6(32'h3cb6cbcf),
	.w7(32'h3c2caaf1),
	.w8(32'hbc0af3d3),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9711014),
	.w1(32'h3c44094b),
	.w2(32'h3b71d3cb),
	.w3(32'h3c7a1c2b),
	.w4(32'hbb593b45),
	.w5(32'hbc08569d),
	.w6(32'hbc9e1ed4),
	.w7(32'hbbee9bed),
	.w8(32'hbb7aaf82),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c813d36),
	.w1(32'hbc4148fa),
	.w2(32'hbd315b0c),
	.w3(32'hba89b98e),
	.w4(32'hbc6eb103),
	.w5(32'hbcb6f750),
	.w6(32'h3cd48a65),
	.w7(32'h3cb3d7b9),
	.w8(32'h3d080f69),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3d84e1),
	.w1(32'hbaddf6ea),
	.w2(32'h3bb789f8),
	.w3(32'hbadb1e1a),
	.w4(32'hbb369abe),
	.w5(32'h3b5ea5ae),
	.w6(32'hbb99649a),
	.w7(32'hbb9ce136),
	.w8(32'hbc13ae86),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8cf9e1),
	.w1(32'h3c1766d1),
	.w2(32'hbc048981),
	.w3(32'h3cc7e922),
	.w4(32'h3ca60e32),
	.w5(32'hbc6c92f4),
	.w6(32'h3b1f3f70),
	.w7(32'h3bf64e1d),
	.w8(32'hba741fac),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0e2ba9),
	.w1(32'h3b6ef361),
	.w2(32'hbbfdb817),
	.w3(32'hbc58fe68),
	.w4(32'h3cd446b5),
	.w5(32'hbcb78000),
	.w6(32'h3b95a2eb),
	.w7(32'h3b674212),
	.w8(32'h3c9d7d53),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc68ec50),
	.w1(32'hbc72e703),
	.w2(32'hbba8ae9c),
	.w3(32'hbb7bf71c),
	.w4(32'hbb410790),
	.w5(32'h3c6c8236),
	.w6(32'h3bb8bd8f),
	.w7(32'h3bbd59c0),
	.w8(32'h3c5f3d39),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ccea6ab),
	.w1(32'hbc08a4cb),
	.w2(32'hbcb132de),
	.w3(32'h3c4bbdba),
	.w4(32'hbc7e8b7a),
	.w5(32'hbbba7f6d),
	.w6(32'h3c688645),
	.w7(32'hbca8b843),
	.w8(32'h3b7bb93f),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc81ec6d),
	.w1(32'h3ace2b00),
	.w2(32'h3c51a7d7),
	.w3(32'hbc6fe8d0),
	.w4(32'hbbd7a65a),
	.w5(32'hbb9d5d90),
	.w6(32'hbca14869),
	.w7(32'hbbfb5dcd),
	.w8(32'hbbbc1e78),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc738b10),
	.w1(32'h3bf8a05f),
	.w2(32'h3ca50d06),
	.w3(32'hbcbc222d),
	.w4(32'hbc5ee095),
	.w5(32'hbb88570b),
	.w6(32'hbc969433),
	.w7(32'hbb2a08fa),
	.w8(32'h395421e0),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c92d5b8),
	.w1(32'h3c65b9c2),
	.w2(32'hbb1e9651),
	.w3(32'h3b5361ab),
	.w4(32'h3c3d2105),
	.w5(32'h3bcbc6ea),
	.w6(32'h3b21d5f6),
	.w7(32'h3bc82021),
	.w8(32'h3984c793),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2063ae),
	.w1(32'h3aec76cf),
	.w2(32'hbb97d972),
	.w3(32'h3abbe72d),
	.w4(32'hbb8112b8),
	.w5(32'hbba728f9),
	.w6(32'hbc83e9c4),
	.w7(32'hbc6f15c4),
	.w8(32'h3b1b0776),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae7f2de),
	.w1(32'h3aad9944),
	.w2(32'hbbcc47a0),
	.w3(32'hb98a074d),
	.w4(32'h3a4fb145),
	.w5(32'h3b8c29ac),
	.w6(32'hbbad62f5),
	.w7(32'hba42b310),
	.w8(32'h3c49befe),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd26ef3),
	.w1(32'h3c3ff72c),
	.w2(32'hbc5a8911),
	.w3(32'h3c3fb2a0),
	.w4(32'h3c6419a8),
	.w5(32'h3b24b9f3),
	.w6(32'h3ceb1d50),
	.w7(32'h3cc5e54e),
	.w8(32'hbc1d5863),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b552dbf),
	.w1(32'hbb15a3ce),
	.w2(32'h3ca9e53b),
	.w3(32'h3c7b4256),
	.w4(32'h3c9e9642),
	.w5(32'h3c1fd03b),
	.w6(32'hbb7baf33),
	.w7(32'hbab85ab4),
	.w8(32'hba85c750),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5239a3),
	.w1(32'hbbcbff0a),
	.w2(32'h3bc1f0bd),
	.w3(32'h3c63cc0a),
	.w4(32'h3aa684bb),
	.w5(32'h3ca1eef3),
	.w6(32'h3c364190),
	.w7(32'hbc6f70b8),
	.w8(32'h3b41897e),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9920ca),
	.w1(32'h3a46da49),
	.w2(32'h3c013c17),
	.w3(32'h3cb34f74),
	.w4(32'h3c439332),
	.w5(32'h3c4f4540),
	.w6(32'h3b9cc8cb),
	.w7(32'hba3cb494),
	.w8(32'h3c64ea47),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1e0b4a),
	.w1(32'h39a2a11b),
	.w2(32'h3b6d36dc),
	.w3(32'h3cfc028a),
	.w4(32'h3c985a71),
	.w5(32'hbbb25910),
	.w6(32'h3c7fa13d),
	.w7(32'h3b0425c1),
	.w8(32'hbc41b85e),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d0a482d),
	.w1(32'hbc2eb389),
	.w2(32'hbc972714),
	.w3(32'h3cec8c8d),
	.w4(32'h3ae5a898),
	.w5(32'hbc175663),
	.w6(32'h3bc28876),
	.w7(32'hbc83252f),
	.w8(32'h3ad13a61),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1e9698),
	.w1(32'hbbb9824b),
	.w2(32'hbc212b7e),
	.w3(32'h3b6d4548),
	.w4(32'h3b9d7ac7),
	.w5(32'hbc19a3f6),
	.w6(32'h3b7b5bcc),
	.w7(32'h3bc45568),
	.w8(32'hbc3e4895),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2dba22),
	.w1(32'hba1cf1c0),
	.w2(32'hb9df8fff),
	.w3(32'hbca1c676),
	.w4(32'hbc533b02),
	.w5(32'h3a491111),
	.w6(32'hbc83a3c6),
	.w7(32'hbc1d2138),
	.w8(32'hbbfa61ec),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c194c6e),
	.w1(32'h3af143e5),
	.w2(32'hbc600aa8),
	.w3(32'h3c39c908),
	.w4(32'h3b850fe7),
	.w5(32'h3b45958f),
	.w6(32'hbb151613),
	.w7(32'hbbe87593),
	.w8(32'h3ba341ed),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabd41d6),
	.w1(32'h3906d203),
	.w2(32'hbbfff83e),
	.w3(32'h3bd3d288),
	.w4(32'h3bb759b3),
	.w5(32'hbc32e47f),
	.w6(32'h3bb05c77),
	.w7(32'h3c05972c),
	.w8(32'hbb2c5597),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaef393),
	.w1(32'h3a5da77b),
	.w2(32'hbb4445e9),
	.w3(32'hbb1e7374),
	.w4(32'h3b1451da),
	.w5(32'hbb2b723c),
	.w6(32'hbb8178e1),
	.w7(32'hbb8ac29f),
	.w8(32'h3c1c2c1d),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb22c9a7),
	.w1(32'h3b09a34c),
	.w2(32'h39b89054),
	.w3(32'hbb96774d),
	.w4(32'h3b4c526d),
	.w5(32'h3b9a431b),
	.w6(32'h3c26e791),
	.w7(32'h3c40ab97),
	.w8(32'h3c025865),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395f4dca),
	.w1(32'hbbb70d02),
	.w2(32'hbbafac7e),
	.w3(32'h3c8b09ab),
	.w4(32'h3c518442),
	.w5(32'h3b205b0e),
	.w6(32'h3c41345b),
	.w7(32'h3ba8006c),
	.w8(32'h3b2b68f2),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5c9a3a),
	.w1(32'h3c101bca),
	.w2(32'h3b9054e7),
	.w3(32'hbb8b5a3e),
	.w4(32'h3b654a19),
	.w5(32'hbbef40dc),
	.w6(32'h3b9ed189),
	.w7(32'h3be5aa94),
	.w8(32'hbc308928),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce31c18),
	.w1(32'hbd0e7c0c),
	.w2(32'hbce1e439),
	.w3(32'hbcc72958),
	.w4(32'hbcd6a8c0),
	.w5(32'hbc91aa94),
	.w6(32'hbad450d9),
	.w7(32'h3b839291),
	.w8(32'h3c2913cb),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc0f569),
	.w1(32'hb95f7279),
	.w2(32'hbc9f4aa6),
	.w3(32'h3c1aa0f6),
	.w4(32'h3b452a09),
	.w5(32'h3b20a24f),
	.w6(32'hbc8a37fc),
	.w7(32'hbc9fa90f),
	.w8(32'h3a9c8e35),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb45ffd),
	.w1(32'hbc9bed5a),
	.w2(32'hbccb4c4f),
	.w3(32'h3b16ddc1),
	.w4(32'hbb9dbfe8),
	.w5(32'hbbb82934),
	.w6(32'hbb17eba6),
	.w7(32'h3bd7b5eb),
	.w8(32'h3c0bcd22),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4d2a21),
	.w1(32'h3b374707),
	.w2(32'h3ba42c16),
	.w3(32'h3c343081),
	.w4(32'h3cca47d5),
	.w5(32'hbb6cd9dd),
	.w6(32'h3ba11951),
	.w7(32'h3c2aafaa),
	.w8(32'hbc2be2a9),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be2c120),
	.w1(32'h3b2aa5aa),
	.w2(32'h3bec0fc0),
	.w3(32'hbbafd904),
	.w4(32'hbc106fa0),
	.w5(32'hbb9def98),
	.w6(32'hbc933765),
	.w7(32'hbcabb32c),
	.w8(32'h3b936fe9),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b83681b),
	.w1(32'h3bef081c),
	.w2(32'h3b99568b),
	.w3(32'hbb8bcdf9),
	.w4(32'h3a49e040),
	.w5(32'h3aae30ee),
	.w6(32'h3ba421be),
	.w7(32'h3c0bfbb9),
	.w8(32'hbc0e666e),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c01834e),
	.w1(32'h3c03adb2),
	.w2(32'hbb1a6074),
	.w3(32'h3b74c233),
	.w4(32'h3b87b39f),
	.w5(32'h3ac95439),
	.w6(32'hbc4be8a3),
	.w7(32'hbc4245b0),
	.w8(32'h3b52e4fb),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb41e251),
	.w1(32'hbc0d1168),
	.w2(32'hbb61fd71),
	.w3(32'h3ce26582),
	.w4(32'h3cadf661),
	.w5(32'h3cd42498),
	.w6(32'h3c8a2135),
	.w7(32'h3be8e476),
	.w8(32'h3c7fa2f7),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd72283),
	.w1(32'hbb69c7fb),
	.w2(32'hb9d491ba),
	.w3(32'h3cb28ea5),
	.w4(32'h3c17f605),
	.w5(32'hbb33ff28),
	.w6(32'h3c18f2d3),
	.w7(32'h3b8d11f5),
	.w8(32'hb9c4e84b),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1ac4cc),
	.w1(32'h3c107dc9),
	.w2(32'hba9f476d),
	.w3(32'hbb89a925),
	.w4(32'h3b9025ce),
	.w5(32'hbb01dfa0),
	.w6(32'h3bf40f28),
	.w7(32'h3c2a6f21),
	.w8(32'hbb3753c5),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1ec481),
	.w1(32'hbbd1ec38),
	.w2(32'h3b4aafa9),
	.w3(32'hbbc5b902),
	.w4(32'hba8b5112),
	.w5(32'h3a98ca90),
	.w6(32'hbbbb01e4),
	.w7(32'hbacc595c),
	.w8(32'hbb29ca5a),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b65e280),
	.w1(32'h3acdd33c),
	.w2(32'hbb95de87),
	.w3(32'h3bb9c781),
	.w4(32'h3b71ee6f),
	.w5(32'hbbddfa11),
	.w6(32'h3b62bcb4),
	.w7(32'h3b4ccdfa),
	.w8(32'hbbf7d17c),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5caf1e),
	.w1(32'hbbee89bd),
	.w2(32'hbb0403e7),
	.w3(32'hbca7efad),
	.w4(32'hbcdce908),
	.w5(32'hbb2a8179),
	.w6(32'hbcba60f0),
	.w7(32'hbc89a93a),
	.w8(32'hbbaae3fe),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8b03dc),
	.w1(32'h3b29c0ad),
	.w2(32'hbae50488),
	.w3(32'hba463266),
	.w4(32'h3b464fb4),
	.w5(32'h3abde02c),
	.w6(32'hbb832f4c),
	.w7(32'h3b01704d),
	.w8(32'hbc14c89e),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd021c2a),
	.w1(32'hbcc85b54),
	.w2(32'hbc829ab2),
	.w3(32'hbc9aac94),
	.w4(32'hbce13018),
	.w5(32'h3a3b935c),
	.w6(32'hbc58ac31),
	.w7(32'h3b1cf31f),
	.w8(32'h3ca4e985),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c22fa19),
	.w1(32'hbb41d237),
	.w2(32'h3c4471a7),
	.w3(32'h3b84e107),
	.w4(32'h3ad9c989),
	.w5(32'h3b84013d),
	.w6(32'hbbb9be35),
	.w7(32'hbba35853),
	.w8(32'h3b8b6106),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b01dc38),
	.w1(32'hbb0b3c0a),
	.w2(32'hb9c3db0e),
	.w3(32'hbb4fda76),
	.w4(32'hbbf12944),
	.w5(32'hbbed3f38),
	.w6(32'hbcd4ecbb),
	.w7(32'hbbebde7f),
	.w8(32'hbb99d485),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule