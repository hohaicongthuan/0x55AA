module layer_8_featuremap_0(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5f34ef),
	.w1(32'hba90cbdd),
	.w2(32'h3bd570cb),
	.w3(32'h3c222989),
	.w4(32'h3ac66fe5),
	.w5(32'h3b9b8801),
	.w6(32'h3c4bb3aa),
	.w7(32'hbac45e29),
	.w8(32'h3b494749),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7227ae),
	.w1(32'h3bd6a5b1),
	.w2(32'hbc1b9da5),
	.w3(32'hbb57fc50),
	.w4(32'h3c2b5156),
	.w5(32'hbc3ac910),
	.w6(32'hbb849e38),
	.w7(32'h3c2f6f90),
	.w8(32'hbbfe911b),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc445889),
	.w1(32'h3af5aca9),
	.w2(32'hba0e0f24),
	.w3(32'hbc1114a1),
	.w4(32'h3ac37d4a),
	.w5(32'hbbadb47e),
	.w6(32'hbc0753c1),
	.w7(32'h3b782138),
	.w8(32'hbbafe12f),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0fac9b),
	.w1(32'hbb80a60a),
	.w2(32'h39c84892),
	.w3(32'h38ce493b),
	.w4(32'hbb8cd189),
	.w5(32'hbabfe6ff),
	.w6(32'h3b7332be),
	.w7(32'hbb7dc71a),
	.w8(32'h3acc8047),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b36a3fa),
	.w1(32'h3b4136ed),
	.w2(32'h3b8077fc),
	.w3(32'h3a84b510),
	.w4(32'h3befb1d6),
	.w5(32'h3a7688e0),
	.w6(32'h3b8ef3b5),
	.w7(32'h393da555),
	.w8(32'hb9b0e282),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a709d19),
	.w1(32'hba9b61a3),
	.w2(32'h3c123cb7),
	.w3(32'h3a25a075),
	.w4(32'hbc8f2fc8),
	.w5(32'hbc9f49ef),
	.w6(32'hba5d37f5),
	.w7(32'hbc3a3142),
	.w8(32'hbc6db77e),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8e97b1),
	.w1(32'hbbb765f5),
	.w2(32'h39f93ef0),
	.w3(32'hbc50cd3a),
	.w4(32'hbbb96f08),
	.w5(32'h3be62ed3),
	.w6(32'hbbecac39),
	.w7(32'hbc645813),
	.w8(32'hbc136fe7),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb578c7d),
	.w1(32'hbc8bf169),
	.w2(32'hbd1260ca),
	.w3(32'h3bbb4cf3),
	.w4(32'hbc265d0f),
	.w5(32'hbcc97258),
	.w6(32'hbb68b076),
	.w7(32'hbc30d793),
	.w8(32'hbc158137),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc87fa23),
	.w1(32'h3bfb5703),
	.w2(32'h3a58210a),
	.w3(32'hbcbdd50e),
	.w4(32'h3c041651),
	.w5(32'h3abf425a),
	.w6(32'hbc5e168d),
	.w7(32'h3c489d4b),
	.w8(32'h3c0a457e),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb903d114),
	.w1(32'hbc1b8d87),
	.w2(32'hbcc1ccc2),
	.w3(32'hbad91d9f),
	.w4(32'h3aff7c65),
	.w5(32'hbb5e39f1),
	.w6(32'h3bf4bfea),
	.w7(32'h3b7e21ec),
	.w8(32'hbae8f4d5),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcfb7884),
	.w1(32'h3bb95899),
	.w2(32'hbbab1280),
	.w3(32'hbd0c8b5e),
	.w4(32'h3c12a6bf),
	.w5(32'hbb02625d),
	.w6(32'hbcb1f05f),
	.w7(32'h3c14967b),
	.w8(32'h3c11e0e1),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3d33e5),
	.w1(32'hbb5e7d22),
	.w2(32'hbb977ad5),
	.w3(32'hbbf0e1fa),
	.w4(32'hbbf238ef),
	.w5(32'hbb7aaadd),
	.w6(32'h3b854d3d),
	.w7(32'hbc2eaedf),
	.w8(32'hbbf3285f),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7868b9),
	.w1(32'h3ce5c990),
	.w2(32'h3c606e6b),
	.w3(32'h3c9d1b63),
	.w4(32'h3bd878c5),
	.w5(32'h3d394e6f),
	.w6(32'hbabcd568),
	.w7(32'h3c38af08),
	.w8(32'h3cd95ae6),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb7ce7b),
	.w1(32'h3bea47a6),
	.w2(32'hbc31d664),
	.w3(32'h3b9465ca),
	.w4(32'h3c57b4b7),
	.w5(32'hbc9b5045),
	.w6(32'h3cf757c8),
	.w7(32'h3cfd42d9),
	.w8(32'h3c26e7b6),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba548e3),
	.w1(32'hbb08dd19),
	.w2(32'h3ac4a6ac),
	.w3(32'hbca8cc72),
	.w4(32'hbb807015),
	.w5(32'h3ba7fe16),
	.w6(32'h3a11e2c2),
	.w7(32'hbc2694b4),
	.w8(32'hbbf6f5ba),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4ac0c6),
	.w1(32'h3957415f),
	.w2(32'h3bbb841b),
	.w3(32'h3bf4990a),
	.w4(32'h3b809076),
	.w5(32'hbb0c2e80),
	.w6(32'hbb41c988),
	.w7(32'h3c06890e),
	.w8(32'h3bdfc5e8),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bac7706),
	.w1(32'hbc2d7372),
	.w2(32'hbce77a96),
	.w3(32'hbbb99004),
	.w4(32'hbca20716),
	.w5(32'hbcf2da32),
	.w6(32'h3bf56b44),
	.w7(32'hbc42fb6f),
	.w8(32'hbce768e7),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0afc75),
	.w1(32'h3b88e1e1),
	.w2(32'h3b2b57d5),
	.w3(32'h3c054a24),
	.w4(32'h3bc9210c),
	.w5(32'h3aac9406),
	.w6(32'hbb616fbb),
	.w7(32'h3c0b0118),
	.w8(32'h3bc8a593),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99977d9),
	.w1(32'hbbdffd13),
	.w2(32'h3b040c05),
	.w3(32'hbb87e1e2),
	.w4(32'hbb948782),
	.w5(32'h3ca2fb28),
	.w6(32'h3ad05e51),
	.w7(32'hbca0a6da),
	.w8(32'hbbaf427d),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d3b6ae6),
	.w1(32'hbb71b1f2),
	.w2(32'hb919f713),
	.w3(32'h3d3a8fc6),
	.w4(32'hbb37a268),
	.w5(32'h3c1743bf),
	.w6(32'h3cd46e89),
	.w7(32'hbc0b0dbe),
	.w8(32'hbb5bee3d),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6d5607),
	.w1(32'h3be63df4),
	.w2(32'hbc0a0eb1),
	.w3(32'h3c0d049d),
	.w4(32'h3c6b55c9),
	.w5(32'hbc327a67),
	.w6(32'h3ad9aed9),
	.w7(32'h3cce17b3),
	.w8(32'h3c463df6),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba0ab15),
	.w1(32'hbb96b0be),
	.w2(32'h3c45c998),
	.w3(32'hbc128187),
	.w4(32'h3b1b888d),
	.w5(32'hbc1ac0f9),
	.w6(32'h3bca0dba),
	.w7(32'h3c1eae8f),
	.w8(32'hbcaf8b73),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4083b9),
	.w1(32'hbc2bfeda),
	.w2(32'h3be71957),
	.w3(32'hbcbed658),
	.w4(32'h3b8765e0),
	.w5(32'hbb4eca37),
	.w6(32'hbcd50e9a),
	.w7(32'hbba220ad),
	.w8(32'hbca314c4),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbf65ee),
	.w1(32'h3a73c556),
	.w2(32'h3c2f7f3a),
	.w3(32'h3cb740c0),
	.w4(32'hbb547c90),
	.w5(32'h3bdf6220),
	.w6(32'hbb80e670),
	.w7(32'hbc54ea72),
	.w8(32'hbc4fdb53),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3e0c0d),
	.w1(32'h3c81a49d),
	.w2(32'h3c2abe28),
	.w3(32'h3c12871b),
	.w4(32'h3c9e5e21),
	.w5(32'h3bc8e0dd),
	.w6(32'hbc0b24c1),
	.w7(32'h3bd4bd9f),
	.w8(32'h3b3583e9),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b60111d),
	.w1(32'hbaeda015),
	.w2(32'h3c195105),
	.w3(32'h3c0e0cdb),
	.w4(32'hbc6a1c60),
	.w5(32'hbc191862),
	.w6(32'h3c1e6609),
	.w7(32'hbc08b85b),
	.w8(32'hbc81cf33),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca3d9f5),
	.w1(32'h3be798ff),
	.w2(32'hbc178a3a),
	.w3(32'h3c902611),
	.w4(32'h3c4419f9),
	.w5(32'hbc349f59),
	.w6(32'h38c30268),
	.w7(32'h3c590a94),
	.w8(32'hbba57d0a),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa160ea),
	.w1(32'h39807678),
	.w2(32'h3708c7c3),
	.w3(32'hbb262f20),
	.w4(32'hbb167aab),
	.w5(32'hbbff87a0),
	.w6(32'h3b44f758),
	.w7(32'h3bf617a7),
	.w8(32'hbbe3d109),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac72fcb),
	.w1(32'h3ba613ae),
	.w2(32'h3bc312c3),
	.w3(32'h3c181709),
	.w4(32'hbc221d15),
	.w5(32'hbb8ead1c),
	.w6(32'h3b180c2e),
	.w7(32'hbbf34ca1),
	.w8(32'h3acfcfa8),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc243c1),
	.w1(32'hbba2ba25),
	.w2(32'hbc25951f),
	.w3(32'h3b8221d2),
	.w4(32'hbb623556),
	.w5(32'hbb8af5c3),
	.w6(32'h3c2119c4),
	.w7(32'hbc03a55a),
	.w8(32'hbc180c45),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf6b209),
	.w1(32'h3b992f78),
	.w2(32'h3c2e08c6),
	.w3(32'hbb200ae6),
	.w4(32'h3b661cc8),
	.w5(32'h3a317e19),
	.w6(32'hbb914f14),
	.w7(32'hbacab03d),
	.w8(32'h3b7c1f20),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c009684),
	.w1(32'hbbc6760f),
	.w2(32'hbb5c6d61),
	.w3(32'h3b15dada),
	.w4(32'hbb51c8e3),
	.w5(32'hbb2b2d50),
	.w6(32'h3c0afd4e),
	.w7(32'hbc0dacf4),
	.w8(32'hbc1594ae),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af796dc),
	.w1(32'h3b992a13),
	.w2(32'h3a7d3dad),
	.w3(32'hba99ce96),
	.w4(32'h3baf6a7e),
	.w5(32'h3b05425f),
	.w6(32'hbc01362e),
	.w7(32'h3b9e245e),
	.w8(32'h3ab6cdda),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b54274d),
	.w1(32'hbc957f13),
	.w2(32'h3b9cc165),
	.w3(32'h3ae74cd8),
	.w4(32'hbcc5ef3b),
	.w5(32'hbc858e0f),
	.w6(32'h3b4d6c4b),
	.w7(32'hbc614215),
	.w8(32'hbd0e9c57),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfaa815),
	.w1(32'h391cf2c0),
	.w2(32'hbae5f15c),
	.w3(32'h3caedb66),
	.w4(32'hba7cac6e),
	.w5(32'hbba84e9f),
	.w6(32'hbba1ca81),
	.w7(32'h3b69ccfe),
	.w8(32'h39ffc100),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bf13be),
	.w1(32'hb939d05a),
	.w2(32'h3c303bcf),
	.w3(32'hbb8cad0a),
	.w4(32'hbbb4af67),
	.w5(32'h3c0100fb),
	.w6(32'h3a9678b1),
	.w7(32'hbbff2420),
	.w8(32'hbb451796),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8be547),
	.w1(32'h3bd6786a),
	.w2(32'h3ca0f83a),
	.w3(32'h39131551),
	.w4(32'h3c704ec8),
	.w5(32'h3d29d177),
	.w6(32'h3ae50662),
	.w7(32'hbb85c2d9),
	.w8(32'h3c638266),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcab18c4),
	.w1(32'hbc0c53e7),
	.w2(32'hbceba996),
	.w3(32'hb89783e1),
	.w4(32'h3bfcb3eb),
	.w5(32'hbc584c36),
	.w6(32'hbad42115),
	.w7(32'hbb377b1f),
	.w8(32'hbc9ec891),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb0cc5e),
	.w1(32'h3b7b380d),
	.w2(32'h3c1affdf),
	.w3(32'hbd32c1a3),
	.w4(32'h3b7db317),
	.w5(32'h3b8df572),
	.w6(32'hbcdabc9e),
	.w7(32'hbc207dca),
	.w8(32'hbc419bb8),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c60e82c),
	.w1(32'h3b0c5848),
	.w2(32'h3c29505b),
	.w3(32'h3cb04851),
	.w4(32'hbc350211),
	.w5(32'h3c308ba5),
	.w6(32'hba5a9da2),
	.w7(32'hbbc845fb),
	.w8(32'h3b7389d4),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c637d21),
	.w1(32'hbac3c80e),
	.w2(32'hbb25c15c),
	.w3(32'h3c78302a),
	.w4(32'hbc158b59),
	.w5(32'h3b8d93a9),
	.w6(32'h3c2f91ac),
	.w7(32'hbca3705f),
	.w8(32'hbc56b59c),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2f3e9a),
	.w1(32'hbaaaa8ac),
	.w2(32'hbc5fdbbb),
	.w3(32'h3bd7dc5e),
	.w4(32'h3b3681d9),
	.w5(32'hbc81b1fa),
	.w6(32'hbc3347ca),
	.w7(32'h3c554779),
	.w8(32'hb9955cd7),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1ace03),
	.w1(32'h3b9de373),
	.w2(32'h3b0982fb),
	.w3(32'hbc03ff54),
	.w4(32'h3b70122e),
	.w5(32'hb9b78346),
	.w6(32'h3a4aa10d),
	.w7(32'h3bd53880),
	.w8(32'h3b120010),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8e5f2d),
	.w1(32'hbc0f453b),
	.w2(32'h3be7247a),
	.w3(32'h3aae8704),
	.w4(32'hbc58b191),
	.w5(32'hbc076028),
	.w6(32'h3b71185e),
	.w7(32'h3bb34c78),
	.w8(32'hbc335f36),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c68c3b2),
	.w1(32'hbc4b8b7f),
	.w2(32'hbcbe8a65),
	.w3(32'h3c075fa3),
	.w4(32'hba93b1f8),
	.w5(32'h3bc6e7e7),
	.w6(32'hbb152bdd),
	.w7(32'h3bb94750),
	.w8(32'h3ce9f714),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf93aa0),
	.w1(32'hbc88840b),
	.w2(32'h3be9fe8d),
	.w3(32'h3c44f568),
	.w4(32'hbc684b6e),
	.w5(32'h3caf580c),
	.w6(32'h3d2ce2fa),
	.w7(32'hbca6887f),
	.w8(32'h3ca6fad3),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca72062),
	.w1(32'hbb9886b9),
	.w2(32'hbca81dfa),
	.w3(32'h3d1e50f5),
	.w4(32'hbc53a72e),
	.w5(32'hbcd6a264),
	.w6(32'h3d37da50),
	.w7(32'hbc68f890),
	.w8(32'hbcd6076c),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4ca064),
	.w1(32'hbc593143),
	.w2(32'h3c229272),
	.w3(32'hbba9dc3e),
	.w4(32'hbc4a7a5c),
	.w5(32'hbc3aa28c),
	.w6(32'hbc4a13e7),
	.w7(32'hbb1e46a1),
	.w8(32'hbc9d550f),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca554f0),
	.w1(32'hbb9d5979),
	.w2(32'h3baa274d),
	.w3(32'h3cb2cf06),
	.w4(32'hbc24465e),
	.w5(32'h3bc6d74c),
	.w6(32'h3b9a428d),
	.w7(32'hbc770714),
	.w8(32'hbc14d441),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6f3b0a),
	.w1(32'hb9936f18),
	.w2(32'hbc182c2d),
	.w3(32'h3912cc24),
	.w4(32'hbb98119a),
	.w5(32'hbc2730f9),
	.w6(32'hbbeebcde),
	.w7(32'hbbce47f4),
	.w8(32'hbc1fd623),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbee1caf),
	.w1(32'hbbcda4c5),
	.w2(32'hbb4736f2),
	.w3(32'hba2b58a7),
	.w4(32'hbc202961),
	.w5(32'h3bf194d8),
	.w6(32'hbb3d5e10),
	.w7(32'hbc1d5812),
	.w8(32'h37eae741),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6c5252),
	.w1(32'h3b727aff),
	.w2(32'h3af37dbf),
	.w3(32'h3c165889),
	.w4(32'hb8c9ecad),
	.w5(32'h38026305),
	.w6(32'h3b41a83a),
	.w7(32'h3b5b8617),
	.w8(32'h3b735424),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c006f4a),
	.w1(32'h3c8deaa8),
	.w2(32'h3c7a19c2),
	.w3(32'h3ba1ec3b),
	.w4(32'h3c3e8c0d),
	.w5(32'h3c86ef0a),
	.w6(32'h3bd61139),
	.w7(32'h3c093e16),
	.w8(32'h3c9881b9),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c161f82),
	.w1(32'h3b6238b4),
	.w2(32'hbb6e2abc),
	.w3(32'h3cf7dbce),
	.w4(32'hbc3141c2),
	.w5(32'hbcfb7e3d),
	.w6(32'h3c9f8490),
	.w7(32'hbc30b418),
	.w8(32'hbc6b15a1),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b62dd7e),
	.w1(32'hbc48eafc),
	.w2(32'h3cac3c2b),
	.w3(32'h3be17e61),
	.w4(32'hbd20c90a),
	.w5(32'h3c8483d3),
	.w6(32'h3b54f137),
	.w7(32'hbd3a312a),
	.w8(32'hbcae8914),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c420cbc),
	.w1(32'h3b2e3cc4),
	.w2(32'h39c73262),
	.w3(32'h3be71c38),
	.w4(32'h3b73a8f4),
	.w5(32'hba3d7001),
	.w6(32'hbc14b272),
	.w7(32'h3c0910fc),
	.w8(32'h3baa9543),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3b599d),
	.w1(32'h3aff7a73),
	.w2(32'h3c7be270),
	.w3(32'hba901c47),
	.w4(32'hbbaba1a3),
	.w5(32'h3ca1b863),
	.w6(32'h3b4a9e41),
	.w7(32'hbaf6a188),
	.w8(32'h3c51ac79),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8c584d),
	.w1(32'hbac6e80a),
	.w2(32'hbc294ce0),
	.w3(32'h3c998944),
	.w4(32'hbc520be9),
	.w5(32'hbbbfd8ef),
	.w6(32'h3c82653a),
	.w7(32'hbbe2a960),
	.w8(32'hbbbc3cd6),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbabdd10),
	.w1(32'h3ba586e5),
	.w2(32'h3bb7bc52),
	.w3(32'hba9d7268),
	.w4(32'hba4ebc71),
	.w5(32'h3946f74d),
	.w6(32'hbba7d73b),
	.w7(32'hbb3812ec),
	.w8(32'hbb9ede48),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be164c7),
	.w1(32'h3c293ced),
	.w2(32'h3c855aa1),
	.w3(32'h3a8242ca),
	.w4(32'h3bc1ae7e),
	.w5(32'h3ce82168),
	.w6(32'hbb4dbde1),
	.w7(32'hbac4fd6b),
	.w8(32'h3ba52826),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabbb7f8),
	.w1(32'h3aa5cecb),
	.w2(32'hbb963c07),
	.w3(32'h3c5cdb40),
	.w4(32'h3c39f5d1),
	.w5(32'hbbc53f23),
	.w6(32'h3ca0dea1),
	.w7(32'h3cc746d0),
	.w8(32'h3c84f0bd),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7bced5),
	.w1(32'hbca02517),
	.w2(32'hbc16f40c),
	.w3(32'hbc1523cf),
	.w4(32'hbc83f165),
	.w5(32'hbc3e167c),
	.w6(32'h3cbec3ef),
	.w7(32'hbc9b89cf),
	.w8(32'hbc3d8a62),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acc17d3),
	.w1(32'h3b1e9a69),
	.w2(32'h3a851e64),
	.w3(32'h3ca2dd62),
	.w4(32'h3bb15c84),
	.w5(32'h3b6532cb),
	.w6(32'h3c713d76),
	.w7(32'h3c08c319),
	.w8(32'h3c0f915d),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3bab13),
	.w1(32'hbb282dba),
	.w2(32'hba1e4586),
	.w3(32'hbb10514f),
	.w4(32'hbba0f7a3),
	.w5(32'hbaf525dc),
	.w6(32'h3b74e9ea),
	.w7(32'h3a894643),
	.w8(32'hbc328dd9),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd4d28b),
	.w1(32'h3b1d56a6),
	.w2(32'h3b9135d7),
	.w3(32'h3959ac26),
	.w4(32'h3b74e36c),
	.w5(32'h3a809780),
	.w6(32'h3bd17bda),
	.w7(32'h3b93a569),
	.w8(32'h3b81327f),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b68c62b),
	.w1(32'h3a7df6d6),
	.w2(32'hbc608f9e),
	.w3(32'hbbd054f5),
	.w4(32'hba9fd30e),
	.w5(32'hbc5f8c5d),
	.w6(32'hbb660572),
	.w7(32'h3b975900),
	.w8(32'hbb812325),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc12c43a),
	.w1(32'h3bba2f46),
	.w2(32'hbc0b6a6b),
	.w3(32'hbc1173c9),
	.w4(32'h3c1858e8),
	.w5(32'hbc3c673f),
	.w6(32'hba6c2672),
	.w7(32'h3ca1523e),
	.w8(32'h3be3f019),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc59badf),
	.w1(32'h3b9eaf62),
	.w2(32'hbc4b3b02),
	.w3(32'hbca0545f),
	.w4(32'h3ba8a14d),
	.w5(32'hbc88ffd6),
	.w6(32'hbb76abb0),
	.w7(32'h3cb4b509),
	.w8(32'h3bcf5aeb),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5cd8ee),
	.w1(32'h39451b4b),
	.w2(32'h3b95beb5),
	.w3(32'hbcb0dc01),
	.w4(32'hb984ff5d),
	.w5(32'hbbd0970c),
	.w6(32'hba511941),
	.w7(32'h3a865387),
	.w8(32'hb9cf8757),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd5b15f),
	.w1(32'hbc8c948c),
	.w2(32'h3ba1cf37),
	.w3(32'hbc4038c7),
	.w4(32'hbcade308),
	.w5(32'h3ba7084c),
	.w6(32'hbb88f018),
	.w7(32'hbc8e6f39),
	.w8(32'hbb891499),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d131ffe),
	.w1(32'h3b8eceb9),
	.w2(32'hba0d4896),
	.w3(32'h3cae14b4),
	.w4(32'h3bb41d7b),
	.w5(32'h3b18c128),
	.w6(32'hbb175814),
	.w7(32'h3ac2a7c0),
	.w8(32'h3b005bbb),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba415be),
	.w1(32'hbc2da154),
	.w2(32'h3c640274),
	.w3(32'hba630895),
	.w4(32'hbc9b6770),
	.w5(32'h3c93a4c1),
	.w6(32'h3b5549ff),
	.w7(32'h3a91dead),
	.w8(32'hb934bbf7),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bef435c),
	.w1(32'hba055557),
	.w2(32'h39df2643),
	.w3(32'h3ce8dd28),
	.w4(32'h3b00ac7b),
	.w5(32'h3a64432d),
	.w6(32'h3cc2c1c5),
	.w7(32'h3b9f8fd9),
	.w8(32'h3b71adb3),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b15bce8),
	.w1(32'hbc09b592),
	.w2(32'h3bebcd6b),
	.w3(32'h399ae5b0),
	.w4(32'hbce49b71),
	.w5(32'hbc4809b5),
	.w6(32'h3b50a796),
	.w7(32'hbd22505a),
	.w8(32'hbd1a7e94),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7aa11b),
	.w1(32'hbc06f960),
	.w2(32'hbb827c9e),
	.w3(32'h3bf4b016),
	.w4(32'hbc065954),
	.w5(32'hbbe5c929),
	.w6(32'hbc9e3657),
	.w7(32'hbc20879a),
	.w8(32'hbbfa5065),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9a6c0e),
	.w1(32'h3c05db20),
	.w2(32'h3c68d73d),
	.w3(32'h3ab4ce52),
	.w4(32'hbbdbc7c6),
	.w5(32'hbbe0206a),
	.w6(32'hbbcaab02),
	.w7(32'hbb6adbd4),
	.w8(32'hbca43357),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c049b6d),
	.w1(32'h3cea4dfa),
	.w2(32'h3d0e7b9f),
	.w3(32'h3c724d82),
	.w4(32'h3c7c2fc8),
	.w5(32'h3d1431c9),
	.w6(32'hbc933517),
	.w7(32'hbc933f17),
	.w8(32'h3c456cb2),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb64ec69),
	.w1(32'hbbc9997f),
	.w2(32'hbae34893),
	.w3(32'h3c6e09a5),
	.w4(32'hbb83ce55),
	.w5(32'h3b70a9f8),
	.w6(32'h3cd1a075),
	.w7(32'hbbdfbcdd),
	.w8(32'hba972b2f),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1597cb),
	.w1(32'hbbaeb37a),
	.w2(32'h3b1f433a),
	.w3(32'h3c3e3ff3),
	.w4(32'hbc18148c),
	.w5(32'hbbc265c5),
	.w6(32'h3adb8928),
	.w7(32'hbc210f41),
	.w8(32'hbc41244c),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b40d852),
	.w1(32'hbc0479df),
	.w2(32'hbb1b17fa),
	.w3(32'h3b21976f),
	.w4(32'hbab0d4ba),
	.w5(32'h3b0d7ba3),
	.w6(32'hbbc7a992),
	.w7(32'hba98acdc),
	.w8(32'hba1a69c9),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be46052),
	.w1(32'hbca388f5),
	.w2(32'hbc83334c),
	.w3(32'h3c70b38e),
	.w4(32'hbc646232),
	.w5(32'hbd0030ac),
	.w6(32'hba559496),
	.w7(32'hbc92bdb1),
	.w8(32'hbce2ed94),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5223cc),
	.w1(32'hbb5b62e3),
	.w2(32'hbac99483),
	.w3(32'hbb9ac4a1),
	.w4(32'hbb935d5b),
	.w5(32'hbae8b100),
	.w6(32'hbc8e8517),
	.w7(32'hbbbd1762),
	.w8(32'hbba37a1a),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcf9a34),
	.w1(32'hbc816851),
	.w2(32'hbc5b2e91),
	.w3(32'h3b9daa83),
	.w4(32'hbbd49ce6),
	.w5(32'hbca4d9f9),
	.w6(32'hbb5953a1),
	.w7(32'h3c463b1f),
	.w8(32'hbbda3325),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bef609f),
	.w1(32'h3b9c0ba0),
	.w2(32'h3b86c1cf),
	.w3(32'hb9d95c72),
	.w4(32'h3b6dc6e3),
	.w5(32'h3b079e8c),
	.w6(32'hbbbc17fd),
	.w7(32'h3be46249),
	.w8(32'h3ba07353),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fdd498),
	.w1(32'hbbad7e3c),
	.w2(32'hbb8d6f78),
	.w3(32'h3a921652),
	.w4(32'hbb01b057),
	.w5(32'hba5781ad),
	.w6(32'h3baf2564),
	.w7(32'hbb4f3c01),
	.w8(32'hbbbeafba),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5446cd),
	.w1(32'hbcbf2568),
	.w2(32'hbcb9c208),
	.w3(32'h3b977243),
	.w4(32'hbbbbf91e),
	.w5(32'hbcaa51bd),
	.w6(32'hbb9ada2c),
	.w7(32'hbb7632b3),
	.w8(32'hb93ef349),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcee1d92),
	.w1(32'h3c06c602),
	.w2(32'h3c4499f9),
	.w3(32'hbc982bbb),
	.w4(32'hb908e167),
	.w5(32'h3b904e5d),
	.w6(32'h3b834779),
	.w7(32'hbb933594),
	.w8(32'hbbe58a9f),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c267ef5),
	.w1(32'h3b0b8651),
	.w2(32'hbb7297ad),
	.w3(32'h3c880068),
	.w4(32'h3b8bc2e0),
	.w5(32'hba830e39),
	.w6(32'h3c0c2323),
	.w7(32'h3b848174),
	.w8(32'h3b21b201),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbf571e),
	.w1(32'hbb4cb85f),
	.w2(32'h3c4f2dc2),
	.w3(32'hbae1d267),
	.w4(32'h3bab7a2f),
	.w5(32'h3ab96f39),
	.w6(32'h3af74c14),
	.w7(32'h39d64910),
	.w8(32'hbc441e83),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbd1f96),
	.w1(32'hbb120484),
	.w2(32'hbb5e9e70),
	.w3(32'h3bc87a47),
	.w4(32'hbb806619),
	.w5(32'hbc25f4ce),
	.w6(32'hbc727c95),
	.w7(32'h3b2ef4c2),
	.w8(32'hba95cf12),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb96d5fc),
	.w1(32'h3b6a19f5),
	.w2(32'hbb310547),
	.w3(32'hbbb38ef7),
	.w4(32'h3be25ae6),
	.w5(32'h3a866c54),
	.w6(32'h3bc91f12),
	.w7(32'h3c0a087d),
	.w8(32'h3b06728d),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbf6d2e),
	.w1(32'hbbd38f6f),
	.w2(32'h3c0279cf),
	.w3(32'h3bff8cae),
	.w4(32'hbb0e0eed),
	.w5(32'h3c951f4b),
	.w6(32'h3bc27dfd),
	.w7(32'hbbed199c),
	.w8(32'h3c01af35),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5a0925),
	.w1(32'hbbf55d99),
	.w2(32'h3a71d949),
	.w3(32'h3cb15494),
	.w4(32'hbc937e41),
	.w5(32'hbc5ad0d1),
	.w6(32'h3c4e80ec),
	.w7(32'hbc5325c9),
	.w8(32'hbccbb524),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7796f0),
	.w1(32'h3aa614dc),
	.w2(32'hba074bbe),
	.w3(32'h3a73cdf4),
	.w4(32'h3a102f1c),
	.w5(32'h3b635296),
	.w6(32'hbc43da36),
	.w7(32'hbb08ba42),
	.w8(32'hbb0755ec),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a610255),
	.w1(32'hbb83f21a),
	.w2(32'h3bf8d017),
	.w3(32'h3b32da12),
	.w4(32'hbbbecf4d),
	.w5(32'hbbdd3832),
	.w6(32'hbb09c2d6),
	.w7(32'hbbee68c9),
	.w8(32'hbc1c46c9),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1703c1),
	.w1(32'h3b0f665c),
	.w2(32'h3a5d26e0),
	.w3(32'h3be127d8),
	.w4(32'h38b1342e),
	.w5(32'h3a5e78de),
	.w6(32'hbc70ba47),
	.w7(32'h3b37fb04),
	.w8(32'h3ac0e0b0),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b59d9de),
	.w1(32'hbb326a54),
	.w2(32'hbb0fac2a),
	.w3(32'h3a943c95),
	.w4(32'hbaf07c7a),
	.w5(32'hba3b53d5),
	.w6(32'h3b8b297c),
	.w7(32'hbb1dac2b),
	.w8(32'h3a5316f7),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3dc377),
	.w1(32'h3c15cf3f),
	.w2(32'h3c21af35),
	.w3(32'hb9e69fd8),
	.w4(32'h3c7561f5),
	.w5(32'h3cad842b),
	.w6(32'h3a8400ba),
	.w7(32'hbb147256),
	.w8(32'h3b8a08bd),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbacca1),
	.w1(32'hba6ac7ef),
	.w2(32'hbb3d0d89),
	.w3(32'h3c5b6201),
	.w4(32'hba9f0c0f),
	.w5(32'h3947b810),
	.w6(32'h3b945cf9),
	.w7(32'hba3c82c9),
	.w8(32'hbaeed437),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba82ea35),
	.w1(32'h3abe1b30),
	.w2(32'h3adb42f4),
	.w3(32'h3a4109bd),
	.w4(32'hbb1e0788),
	.w5(32'hbb70f480),
	.w6(32'hba65008e),
	.w7(32'hbc08063e),
	.w8(32'hbc23597f),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf065b6),
	.w1(32'hbc5165f2),
	.w2(32'hbb270142),
	.w3(32'h3af08e1b),
	.w4(32'hbc9c3e7b),
	.w5(32'hbca69494),
	.w6(32'hbbd1e07c),
	.w7(32'hbc85f7f5),
	.w8(32'hbca2c983),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a15aa14),
	.w1(32'hbc125768),
	.w2(32'h3b7a1a17),
	.w3(32'hbc4220fd),
	.w4(32'hbcc8f80d),
	.w5(32'h3c225f91),
	.w6(32'hbc5d2a2d),
	.w7(32'hbcbac9b8),
	.w8(32'hbc59515c),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cac259a),
	.w1(32'hbbed20f7),
	.w2(32'h3bda9c0b),
	.w3(32'h3c1be273),
	.w4(32'hbc74fb95),
	.w5(32'h375c1c39),
	.w6(32'h3b8a8cec),
	.w7(32'hbc8d6152),
	.w8(32'hbc268ecd),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c264988),
	.w1(32'hbb74775a),
	.w2(32'h3b9ed6b8),
	.w3(32'h3c729bb2),
	.w4(32'hbbdf04a3),
	.w5(32'h3aaa59ce),
	.w6(32'h3be07cf5),
	.w7(32'hbbe23885),
	.w8(32'hbc1d4c78),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdfbd1b),
	.w1(32'hb9b8ea82),
	.w2(32'hbb4de54f),
	.w3(32'hbb3ab84c),
	.w4(32'hbb59a8bf),
	.w5(32'h3bdf689d),
	.w6(32'hbc00df4b),
	.w7(32'hbc6ec5ad),
	.w8(32'hbc08c996),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc17b31),
	.w1(32'h398d0a6e),
	.w2(32'h3b0ce5b1),
	.w3(32'h3c44b7f4),
	.w4(32'h3b657f88),
	.w5(32'h3b987156),
	.w6(32'h3b7a4c94),
	.w7(32'h3b6e8a67),
	.w8(32'h3b8cf8b0),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be4b33a),
	.w1(32'h3b2c73b9),
	.w2(32'h3b782db3),
	.w3(32'h3bfeee87),
	.w4(32'h3b03c500),
	.w5(32'h3b8af80f),
	.w6(32'h3b91170c),
	.w7(32'h39e90fd6),
	.w8(32'h3b46620b),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabed2ef),
	.w1(32'h3a8420ee),
	.w2(32'hbc1ae9af),
	.w3(32'h3aef3abe),
	.w4(32'hbbdf25d2),
	.w5(32'h3bd4667b),
	.w6(32'h3b3b7019),
	.w7(32'hbbed5bbe),
	.w8(32'hbbc3c483),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf247ac),
	.w1(32'h3b0587e4),
	.w2(32'hbbe497e7),
	.w3(32'h3bf63466),
	.w4(32'h3bcea8f9),
	.w5(32'h3c07611e),
	.w6(32'h3b049547),
	.w7(32'h3a0333aa),
	.w8(32'hbb322e60),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4923c5),
	.w1(32'h3c5f1160),
	.w2(32'h3c216eed),
	.w3(32'h3aedfe70),
	.w4(32'h3a9aac30),
	.w5(32'h3bcba55c),
	.w6(32'hbbf900b6),
	.w7(32'h3bfeeccb),
	.w8(32'h3ac7f6b4),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7a8d9f),
	.w1(32'h3a60bf1b),
	.w2(32'h3ba30368),
	.w3(32'h3bbfb41d),
	.w4(32'hbc1e3419),
	.w5(32'hbb8321fe),
	.w6(32'hbc4a8484),
	.w7(32'hbc5e52fa),
	.w8(32'hbce0b2d6),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5470d7),
	.w1(32'h3c11184e),
	.w2(32'h3b6c8cf0),
	.w3(32'hba21c5e8),
	.w4(32'hbb122f1b),
	.w5(32'h3c20f963),
	.w6(32'hbcbfe750),
	.w7(32'hbbad58c6),
	.w8(32'h3a3f4a99),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbcb528),
	.w1(32'h3a406eea),
	.w2(32'h3a6a536e),
	.w3(32'h3c20e4b0),
	.w4(32'hbb9c06b9),
	.w5(32'hbbd08506),
	.w6(32'h3aa793aa),
	.w7(32'hbbb4a8f5),
	.w8(32'hbc103b5f),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a99eb1c),
	.w1(32'hbbc26242),
	.w2(32'hbbb172f8),
	.w3(32'hba3bec20),
	.w4(32'hb966f97c),
	.w5(32'hbbdc8f52),
	.w6(32'hbb469f80),
	.w7(32'hbb2faac1),
	.w8(32'hb7ffb6bd),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb340c24),
	.w1(32'h3b1f35dd),
	.w2(32'h3bbfa6d7),
	.w3(32'h3ab4d977),
	.w4(32'hbaa78e5b),
	.w5(32'hbbae7923),
	.w6(32'hbb94e260),
	.w7(32'hbb2f040d),
	.w8(32'hbbb0c6e3),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5255e5),
	.w1(32'h39e888ee),
	.w2(32'h3b9ba195),
	.w3(32'h3ac456c0),
	.w4(32'h3947b9c2),
	.w5(32'h3b84712e),
	.w6(32'hbb725be5),
	.w7(32'hbace600b),
	.w8(32'h3af96091),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b39e839),
	.w1(32'hbbb345ef),
	.w2(32'h3c06dd17),
	.w3(32'h3b54a7af),
	.w4(32'hbb7e6fd9),
	.w5(32'hbb45eb1e),
	.w6(32'h3af7a189),
	.w7(32'hbb8cb7d1),
	.w8(32'hbb2fb8e1),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d08e60c),
	.w1(32'h3bfd27ee),
	.w2(32'h3b3f82a3),
	.w3(32'h3cb22348),
	.w4(32'hbb8a21f4),
	.w5(32'hbc3e0ac0),
	.w6(32'h3c25022f),
	.w7(32'hbc25a007),
	.w8(32'hbc17f894),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c49c23e),
	.w1(32'h3cfcf8a2),
	.w2(32'h3cef89eb),
	.w3(32'hbb05dca6),
	.w4(32'h3ca15703),
	.w5(32'h3d113ad8),
	.w6(32'h3a812eac),
	.w7(32'hbc4b5214),
	.w8(32'h3c9963a9),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3caabb7f),
	.w1(32'hbb1573bf),
	.w2(32'hb9c77b2d),
	.w3(32'h3d0d0d50),
	.w4(32'hbb903985),
	.w5(32'hbaae444c),
	.w6(32'h3cbe902d),
	.w7(32'hbbb0daec),
	.w8(32'hbb9b4eae),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd8b880),
	.w1(32'hbb8d4ed6),
	.w2(32'h3b71722f),
	.w3(32'h3baed831),
	.w4(32'hbc5367e2),
	.w5(32'hbc08dfdc),
	.w6(32'hbaa678ee),
	.w7(32'hbc7c108b),
	.w8(32'hbca074d9),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b285306),
	.w1(32'hbc2e7490),
	.w2(32'h3b676ebf),
	.w3(32'hbb568c96),
	.w4(32'hbc8404b8),
	.w5(32'hbba971e8),
	.w6(32'hbc47385c),
	.w7(32'hbc1d4ecc),
	.w8(32'hbbaa1fc2),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9e33fd),
	.w1(32'hba864137),
	.w2(32'h3af31134),
	.w3(32'h3bfd0c8b),
	.w4(32'hbba4eb8a),
	.w5(32'hba9c8e55),
	.w6(32'hb92f9591),
	.w7(32'hbb4e4a9e),
	.w8(32'hbb02e363),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4f4459),
	.w1(32'hbc03a3f6),
	.w2(32'h3d188816),
	.w3(32'h3b9b5dcf),
	.w4(32'hbd1f56df),
	.w5(32'hbcae5c00),
	.w6(32'hb8108eea),
	.w7(32'hbd5ab4f2),
	.w8(32'hbd48edf1),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d85b191),
	.w1(32'hbaffd275),
	.w2(32'hbbcfd7de),
	.w3(32'h3d168e4d),
	.w4(32'h3b1f08e6),
	.w5(32'h3aaad143),
	.w6(32'hbbe593f9),
	.w7(32'h3aec4578),
	.w8(32'hbac97fd5),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1ce443),
	.w1(32'h3b2dae6a),
	.w2(32'h3c56d523),
	.w3(32'h3c48e220),
	.w4(32'hbc94b78d),
	.w5(32'h3c16df35),
	.w6(32'h3b2a649d),
	.w7(32'hbc9a938c),
	.w8(32'hbcbe49ad),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3ba52c),
	.w1(32'hbb443413),
	.w2(32'hbac59090),
	.w3(32'h3c538264),
	.w4(32'hbb35d312),
	.w5(32'hbb08e9df),
	.w6(32'hbbcfb6d9),
	.w7(32'h3a01130e),
	.w8(32'hbaa664ca),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aac0fce),
	.w1(32'hbbfcae51),
	.w2(32'hbc20eb87),
	.w3(32'hb9e06f4f),
	.w4(32'hba07bb6b),
	.w5(32'hbcddd970),
	.w6(32'hba70624b),
	.w7(32'hba8dddf1),
	.w8(32'hbc95f632),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule