module layer_8_featuremap_132(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b13a40d),
	.w1(32'h3c3386e3),
	.w2(32'h3cac2d2f),
	.w3(32'h3b9fc75b),
	.w4(32'h3c6d6df6),
	.w5(32'h3c20c4b1),
	.w6(32'hbaac2e60),
	.w7(32'h3c6870b1),
	.w8(32'hbc2b1de2),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b636cb9),
	.w1(32'h3be7c04d),
	.w2(32'hbb135e01),
	.w3(32'h3b8e5db7),
	.w4(32'h3a8a9fec),
	.w5(32'hbcd0721d),
	.w6(32'hbb9309dc),
	.w7(32'h3bc79166),
	.w8(32'hbc4017bd),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc805376),
	.w1(32'hbc894610),
	.w2(32'h3cafab96),
	.w3(32'hbc9bc7e2),
	.w4(32'h3c57da18),
	.w5(32'hbc2605d5),
	.w6(32'hbc5b3e0a),
	.w7(32'h3c50f74c),
	.w8(32'hbc456f0f),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3e3348),
	.w1(32'hbc1a707f),
	.w2(32'h3b04daa2),
	.w3(32'hbc04ed9f),
	.w4(32'h3a92068c),
	.w5(32'hbcc71bb4),
	.w6(32'hbc85ca35),
	.w7(32'hbbf987bc),
	.w8(32'hbc1953a3),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc80acab),
	.w1(32'hba1c2e9a),
	.w2(32'hbc027c41),
	.w3(32'h3bb96ba4),
	.w4(32'hbc1e465d),
	.w5(32'h3b9f57b8),
	.w6(32'h3bc6a8fc),
	.w7(32'hbc103aa8),
	.w8(32'h3bc4952e),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1ca1fe),
	.w1(32'h3bcebeff),
	.w2(32'hbc6a53b9),
	.w3(32'h3b7c109c),
	.w4(32'hbc260b19),
	.w5(32'hbc63b429),
	.w6(32'hbb983519),
	.w7(32'hbbdd168f),
	.w8(32'h3d0af6b4),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c273cb7),
	.w1(32'h3b9083cc),
	.w2(32'h3c2190cc),
	.w3(32'hb9eee911),
	.w4(32'h3c904982),
	.w5(32'hb92cac18),
	.w6(32'h3c3bb45a),
	.w7(32'h3c5b4600),
	.w8(32'hbc4dc7a0),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba49ef12),
	.w1(32'h3b9549a1),
	.w2(32'h3b99e1ec),
	.w3(32'hbc12758e),
	.w4(32'h3c71914f),
	.w5(32'hbc071b43),
	.w6(32'hbc26da45),
	.w7(32'h3c212263),
	.w8(32'hbc7c0b46),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc230034),
	.w1(32'h38d4423d),
	.w2(32'hbb313fd3),
	.w3(32'hbbb63773),
	.w4(32'hbbd83ba3),
	.w5(32'h3bc2979b),
	.w6(32'hba012766),
	.w7(32'hbac2cb75),
	.w8(32'hbb98127d),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7c77ec),
	.w1(32'h3a4df5f0),
	.w2(32'hbafc2424),
	.w3(32'hbbf2451f),
	.w4(32'hbc93d304),
	.w5(32'hbc311d3f),
	.w6(32'hbc11a3d0),
	.w7(32'h3b88e1b6),
	.w8(32'h3cd70ef1),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9734ea),
	.w1(32'hbbdf5496),
	.w2(32'hbaf82fa2),
	.w3(32'h3b53163e),
	.w4(32'hbb99f250),
	.w5(32'hbba1bde5),
	.w6(32'h3c48da30),
	.w7(32'h3bdb5dc2),
	.w8(32'hbc167dc6),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5c9bcf),
	.w1(32'h3c0f6b79),
	.w2(32'hbb9fa37e),
	.w3(32'h3a63847f),
	.w4(32'h39e662a8),
	.w5(32'hbc3edf12),
	.w6(32'h3bde99b5),
	.w7(32'hbbd82468),
	.w8(32'hbc744412),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5b07c7),
	.w1(32'h3b6f41e7),
	.w2(32'hbab02f6f),
	.w3(32'hbc25e53c),
	.w4(32'h39be6691),
	.w5(32'hbaebfd9e),
	.w6(32'hbbb0154e),
	.w7(32'h3a315839),
	.w8(32'hb9e01210),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7cc804c),
	.w1(32'h3ad410ae),
	.w2(32'hbb4aaa78),
	.w3(32'hba080ff3),
	.w4(32'hbb838bb4),
	.w5(32'hbab55823),
	.w6(32'h39efc841),
	.w7(32'hbb96df65),
	.w8(32'hbb07d57c),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf8115e),
	.w1(32'hbb5713ab),
	.w2(32'hbb47cbc4),
	.w3(32'hbb243f50),
	.w4(32'hbaf6e20b),
	.w5(32'hbad9fe4f),
	.w6(32'hb9d3ff44),
	.w7(32'hbb1c6a98),
	.w8(32'hbb3487ae),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6cb2e5),
	.w1(32'hbb5beca6),
	.w2(32'h39a738dc),
	.w3(32'hbb5b56c7),
	.w4(32'hbb844d84),
	.w5(32'hbb22fd35),
	.w6(32'hbb3dd8c4),
	.w7(32'hba962cf3),
	.w8(32'hbac7849c),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399eccde),
	.w1(32'hbbbbd7e4),
	.w2(32'h3bc8d6e0),
	.w3(32'h3ad9901c),
	.w4(32'h3c17be90),
	.w5(32'h3c949681),
	.w6(32'h3b4287c5),
	.w7(32'h37dcb413),
	.w8(32'h3c7ea0d1),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8bc84c),
	.w1(32'h3b89dac8),
	.w2(32'hbc046da0),
	.w3(32'hb9c7c3c1),
	.w4(32'hbc2af2f1),
	.w5(32'hbb611cd3),
	.w6(32'hbb5f28ce),
	.w7(32'hb8b3bdc9),
	.w8(32'hbbf66fad),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4e33a4),
	.w1(32'hbc20eddb),
	.w2(32'hbb90fcb9),
	.w3(32'hbb8aa042),
	.w4(32'hbbe14842),
	.w5(32'hbc058819),
	.w6(32'h39c6760d),
	.w7(32'hbc109aca),
	.w8(32'hbc8fa712),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3664fd),
	.w1(32'hbb7e7bec),
	.w2(32'hbc2c71fd),
	.w3(32'h37522a0a),
	.w4(32'h3aa5011f),
	.w5(32'hbb91002c),
	.w6(32'hba6d9683),
	.w7(32'hbb8ede02),
	.w8(32'hbb02341c),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2f5dac),
	.w1(32'hbc6a9d33),
	.w2(32'hbb848709),
	.w3(32'h3a58da5f),
	.w4(32'hbb542bd9),
	.w5(32'hbba2cd2f),
	.w6(32'hbbae9e10),
	.w7(32'hb987e604),
	.w8(32'h3c2021d4),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b85d125),
	.w1(32'h3b787713),
	.w2(32'hba8155dd),
	.w3(32'h3bbeaa96),
	.w4(32'h3bbb2429),
	.w5(32'hbb987a2d),
	.w6(32'h3ad80415),
	.w7(32'h3b7c55dc),
	.w8(32'hbb968f77),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8e8945),
	.w1(32'hbbc1c11b),
	.w2(32'hbbc9c2f0),
	.w3(32'hbb789177),
	.w4(32'h3b72461e),
	.w5(32'hbc249236),
	.w6(32'hbb84d3e3),
	.w7(32'hbb63e687),
	.w8(32'hbc83cf02),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd82119),
	.w1(32'h398cc682),
	.w2(32'h3b166b3b),
	.w3(32'hbae87179),
	.w4(32'h3acd35e3),
	.w5(32'h3accc4d5),
	.w6(32'hbb649f0b),
	.w7(32'h3b2d2fd2),
	.w8(32'h3ac4bf70),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadcdd5c),
	.w1(32'hbbf6d401),
	.w2(32'hbbb449ff),
	.w3(32'hbb819db5),
	.w4(32'hbc00c27e),
	.w5(32'hbc01df0d),
	.w6(32'hbb98a728),
	.w7(32'hbc0e353b),
	.w8(32'hbbadaf5d),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb23231c),
	.w1(32'hbb6c481a),
	.w2(32'h38afa2ce),
	.w3(32'h3a239672),
	.w4(32'h3c15ca99),
	.w5(32'hbbfaeeba),
	.w6(32'hba48cfbd),
	.w7(32'hbb7d7a81),
	.w8(32'hbc03d02b),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b926d05),
	.w1(32'hbb085085),
	.w2(32'h3bc56324),
	.w3(32'hbbddcb67),
	.w4(32'hbb1c14a0),
	.w5(32'hb974186e),
	.w6(32'hba8c612a),
	.w7(32'hbbc2b4d1),
	.w8(32'h3ba89d55),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb05071),
	.w1(32'hbccbb1a5),
	.w2(32'hbc4d0ed3),
	.w3(32'h3d00e7d3),
	.w4(32'h3be13622),
	.w5(32'hbc612f22),
	.w6(32'h3cf3c5f5),
	.w7(32'h3c48a1b2),
	.w8(32'hbcfbe00b),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb909176),
	.w1(32'hbb6c74d3),
	.w2(32'hba77bfca),
	.w3(32'h3b80f55e),
	.w4(32'h3af5817c),
	.w5(32'hbbcc6ddb),
	.w6(32'hba1620d1),
	.w7(32'hbb9d3a68),
	.w8(32'hbc12b3eb),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b92ca69),
	.w1(32'h3c4a2a31),
	.w2(32'h3b06d3ae),
	.w3(32'hbb7acff5),
	.w4(32'hbad85ef2),
	.w5(32'hbb61ba5f),
	.w6(32'h39f9a5ec),
	.w7(32'hbb8f63d1),
	.w8(32'h3aacc864),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1828bb),
	.w1(32'h3c047d61),
	.w2(32'hb98c59ff),
	.w3(32'h3b0c1fd1),
	.w4(32'h3896b614),
	.w5(32'hbab695cf),
	.w6(32'h3c488f5a),
	.w7(32'h3a8738ab),
	.w8(32'hb9929f36),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb09a309),
	.w1(32'hbb33f7fd),
	.w2(32'hbabde8d8),
	.w3(32'hbb83a52a),
	.w4(32'hbb135eb7),
	.w5(32'hbb790b1d),
	.w6(32'hbb3d33df),
	.w7(32'hb9eeb471),
	.w8(32'hbbc92268),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3a15ce),
	.w1(32'h3bb7599d),
	.w2(32'h3b4419d8),
	.w3(32'h3b48ad41),
	.w4(32'h3c204383),
	.w5(32'hba5362ba),
	.w6(32'h3b56ae34),
	.w7(32'h3c009be1),
	.w8(32'h3aba8a36),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a83fc44),
	.w1(32'h3b898aa5),
	.w2(32'h3bd4668c),
	.w3(32'hbb3352d2),
	.w4(32'h3b11e794),
	.w5(32'h3c6d34aa),
	.w6(32'hbbe00905),
	.w7(32'h3abbc9be),
	.w8(32'h3c77ad48),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3113fe),
	.w1(32'hba863341),
	.w2(32'h3b371b0e),
	.w3(32'h3b8db051),
	.w4(32'h3bd590f1),
	.w5(32'h3aee4891),
	.w6(32'hbac77f21),
	.w7(32'h3ba694b6),
	.w8(32'h3b256cb8),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b91b467),
	.w1(32'hb9eed9c6),
	.w2(32'hbb0e9184),
	.w3(32'h3b258b38),
	.w4(32'h3af9a046),
	.w5(32'hbbc63821),
	.w6(32'h3b5fa08c),
	.w7(32'h3bc8042c),
	.w8(32'h3b1c2f5b),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9b3db1),
	.w1(32'h3b7f1e17),
	.w2(32'hbbd3639e),
	.w3(32'h3ad8fdd0),
	.w4(32'h3acc1a76),
	.w5(32'hbb2dc793),
	.w6(32'h3b828f54),
	.w7(32'hbbec54b3),
	.w8(32'h37586b3f),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4d2866),
	.w1(32'h3bade28b),
	.w2(32'h3b39eb9d),
	.w3(32'hbba55584),
	.w4(32'h3b9c2fb9),
	.w5(32'hba94210f),
	.w6(32'hbab48557),
	.w7(32'h39e9702b),
	.w8(32'hbb176f68),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb389714),
	.w1(32'hba481262),
	.w2(32'hbad73718),
	.w3(32'h3a4753d2),
	.w4(32'h3b88a9a2),
	.w5(32'h397188cd),
	.w6(32'hbab3a1b9),
	.w7(32'h3a97ad95),
	.w8(32'hbbddffa9),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acd61b0),
	.w1(32'h3be9ff16),
	.w2(32'h3a25fec2),
	.w3(32'hbb8f7922),
	.w4(32'h3979a1a6),
	.w5(32'hbb3c28e7),
	.w6(32'h39b2eee0),
	.w7(32'h3b08c67c),
	.w8(32'hbb29b887),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9346ec),
	.w1(32'hbb4be0bf),
	.w2(32'hbb90924d),
	.w3(32'hbb62ae39),
	.w4(32'hbc736671),
	.w5(32'hbc522b06),
	.w6(32'h3aea6dbd),
	.w7(32'hbc57193b),
	.w8(32'hbc42408d),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4e2a19),
	.w1(32'hbc79059e),
	.w2(32'h3b1401a6),
	.w3(32'hba559e41),
	.w4(32'hbbb9fce3),
	.w5(32'hbb33c3cf),
	.w6(32'hbc131230),
	.w7(32'hbbad33d4),
	.w8(32'h3b30e76b),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2db697),
	.w1(32'hbb366265),
	.w2(32'hb97fbd82),
	.w3(32'h3bda7125),
	.w4(32'h3b990a93),
	.w5(32'hbaf53e5b),
	.w6(32'h3ad3c4e8),
	.w7(32'hbb774e7e),
	.w8(32'hbb91608d),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3c5922),
	.w1(32'h3c79ef34),
	.w2(32'hbb775fc3),
	.w3(32'hbc03d494),
	.w4(32'hbaa59d31),
	.w5(32'hbb297f66),
	.w6(32'hbb637a6c),
	.w7(32'hbaac4cfb),
	.w8(32'hbac2eff1),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a94bbda),
	.w1(32'h3a10e4a8),
	.w2(32'hbb32d908),
	.w3(32'h3a699772),
	.w4(32'hba479bf3),
	.w5(32'hbb99637b),
	.w6(32'h3b67e9c8),
	.w7(32'hbbec28ea),
	.w8(32'hbc1149db),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf3b82e),
	.w1(32'h3bc291be),
	.w2(32'hbb964299),
	.w3(32'hbb8d940c),
	.w4(32'hbacb86b1),
	.w5(32'hbc44c680),
	.w6(32'hbaeeb0e1),
	.w7(32'hbad97f92),
	.w8(32'hbc72ea9c),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb8be84),
	.w1(32'h3c44dcd0),
	.w2(32'hbbd99451),
	.w3(32'h3b46f20f),
	.w4(32'hba6dbcfe),
	.w5(32'hbbb0765e),
	.w6(32'h3ba707b3),
	.w7(32'hbb53a37b),
	.w8(32'hbbff57fa),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b009c16),
	.w1(32'h3a0daa8e),
	.w2(32'h3b1c587a),
	.w3(32'h3b3ec215),
	.w4(32'h3b876abe),
	.w5(32'hbbe8c84d),
	.w6(32'h3b9a5177),
	.w7(32'hbbb1b096),
	.w8(32'hbc053c7f),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be03a1c),
	.w1(32'hba397ed1),
	.w2(32'h3bb49f4a),
	.w3(32'hbc1d07af),
	.w4(32'hbb58c8a2),
	.w5(32'h39f083fd),
	.w6(32'hbb3116f8),
	.w7(32'h3bcf9b40),
	.w8(32'h3af80d09),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae56c34),
	.w1(32'hbb9f4853),
	.w2(32'h3aa33c66),
	.w3(32'h3b5481b0),
	.w4(32'h3a1e6a00),
	.w5(32'h3bbcb05d),
	.w6(32'h3b94ca3c),
	.w7(32'hba7f34f8),
	.w8(32'h3a0a2e68),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b98cfbc),
	.w1(32'h3b936841),
	.w2(32'h3c0f34ff),
	.w3(32'h3b833972),
	.w4(32'h3bde139f),
	.w5(32'h3c251dfb),
	.w6(32'h3c17fd39),
	.w7(32'h3ba3a698),
	.w8(32'h3c23f263),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcc5796),
	.w1(32'hbc20df75),
	.w2(32'hbbb96fe2),
	.w3(32'h3c2222d7),
	.w4(32'h3b723907),
	.w5(32'h3b6523c7),
	.w6(32'h3a300639),
	.w7(32'h3a190b2d),
	.w8(32'h3b330256),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1ee96a),
	.w1(32'h3b701f68),
	.w2(32'hba866e4e),
	.w3(32'h39cc00d2),
	.w4(32'hbc0cd678),
	.w5(32'h3bf2817f),
	.w6(32'hbadb8a73),
	.w7(32'hbb5eeecf),
	.w8(32'h3ab4e920),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba15a465),
	.w1(32'hbb12a42c),
	.w2(32'hbb13140b),
	.w3(32'hb9605ff9),
	.w4(32'hbb773a76),
	.w5(32'hbb862f04),
	.w6(32'hbb88d086),
	.w7(32'hbb18737b),
	.w8(32'hbae47a88),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab53ba7),
	.w1(32'h3aad8c5e),
	.w2(32'hbb44f2ae),
	.w3(32'hb80f38eb),
	.w4(32'hbb8f0ffe),
	.w5(32'hbc049c40),
	.w6(32'h3b02e0b6),
	.w7(32'hbbc25936),
	.w8(32'hbacf3959),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb86f5d88),
	.w1(32'h398c9f1b),
	.w2(32'hbba69d0f),
	.w3(32'h3b8d357a),
	.w4(32'hbb8752a7),
	.w5(32'hbb67d6b3),
	.w6(32'h3b663ce9),
	.w7(32'hbbaeeb12),
	.w8(32'hbbff8063),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b82a852),
	.w1(32'hbb24074d),
	.w2(32'h3c810b3e),
	.w3(32'hbbd04507),
	.w4(32'hbad9a630),
	.w5(32'h3bf15f03),
	.w6(32'hbb85ce44),
	.w7(32'h3c4bac3c),
	.w8(32'h3cb34610),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfb8cac),
	.w1(32'hbb281448),
	.w2(32'h3bf83d38),
	.w3(32'h3c6bce2e),
	.w4(32'hb91e8fbc),
	.w5(32'hbad017c7),
	.w6(32'h3c28d25c),
	.w7(32'h3b780543),
	.w8(32'h3b5d9aa8),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc137b95),
	.w1(32'hbc0b3787),
	.w2(32'hbb368314),
	.w3(32'h3b9313d0),
	.w4(32'hbaf799b3),
	.w5(32'hba04344e),
	.w6(32'h39b3b469),
	.w7(32'hbaf051bc),
	.w8(32'hb9fe703b),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba336d33),
	.w1(32'hb9a61831),
	.w2(32'hbb9903f2),
	.w3(32'hb96458be),
	.w4(32'h3b4f08d5),
	.w5(32'h3b57d7a5),
	.w6(32'hb9df726b),
	.w7(32'h3b90ee66),
	.w8(32'hbbd25cf8),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3783de7d),
	.w1(32'h3abfc3cb),
	.w2(32'h3ba79e67),
	.w3(32'hbc37cbc2),
	.w4(32'h3a84db74),
	.w5(32'h3ae76817),
	.w6(32'hbbdc6aea),
	.w7(32'h3b17dd25),
	.w8(32'h39d9de57),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc232017),
	.w1(32'hbaadfa1b),
	.w2(32'hbabd3e0f),
	.w3(32'h3c049953),
	.w4(32'h3bd62f63),
	.w5(32'h3bf0fa34),
	.w6(32'hbc13bdce),
	.w7(32'h39fbd62a),
	.w8(32'h3bcb90bd),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd09546),
	.w1(32'h3aa0fc71),
	.w2(32'hbc033d62),
	.w3(32'hbba772c7),
	.w4(32'hbc2ca8bb),
	.w5(32'hbc0ca872),
	.w6(32'h3a3ddb06),
	.w7(32'hbc29faa6),
	.w8(32'hbc05fcde),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeeedf0),
	.w1(32'hbc12df87),
	.w2(32'hbb89c3bf),
	.w3(32'hbc2b56a7),
	.w4(32'h3b0937a2),
	.w5(32'hb93ce8bc),
	.w6(32'hbc3fd1dd),
	.w7(32'hba846562),
	.w8(32'hbb66f7ba),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a640022),
	.w1(32'h3b572c5b),
	.w2(32'hbb884e32),
	.w3(32'hba0bf5c8),
	.w4(32'h3b91bf67),
	.w5(32'hbb65c065),
	.w6(32'hbafe7310),
	.w7(32'hbb1503bd),
	.w8(32'hbbfae357),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba9b0cb),
	.w1(32'hba3f1082),
	.w2(32'h3c03f905),
	.w3(32'hbb30562c),
	.w4(32'h3c3a283c),
	.w5(32'h3c796e08),
	.w6(32'hbaf3da2b),
	.w7(32'h3bf3bfe7),
	.w8(32'h3c6a4c51),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c668bf8),
	.w1(32'h3abebe9f),
	.w2(32'hbb9322de),
	.w3(32'hbb2f9a1c),
	.w4(32'hbb3e639f),
	.w5(32'hbbfec564),
	.w6(32'hbb96df0e),
	.w7(32'hbb2d750c),
	.w8(32'hbc48009c),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb06f592),
	.w1(32'h3a386b98),
	.w2(32'hbbce60d7),
	.w3(32'hbaafaf33),
	.w4(32'hbb9b4150),
	.w5(32'hba7916c7),
	.w6(32'h3a847d17),
	.w7(32'hbbc2e504),
	.w8(32'hbb8f47be),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5ff9ee),
	.w1(32'h3beabec7),
	.w2(32'hb93c99ac),
	.w3(32'h386f08e3),
	.w4(32'h38ce4685),
	.w5(32'h3c20a1ad),
	.w6(32'hbc05dc27),
	.w7(32'h3b6582b5),
	.w8(32'hbb9efcf6),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98429af),
	.w1(32'hbbedcdf8),
	.w2(32'h3b740b9c),
	.w3(32'h3c222d42),
	.w4(32'hbb3dae1c),
	.w5(32'h3c28519e),
	.w6(32'h3b945550),
	.w7(32'h38d9fc02),
	.w8(32'h3c78dae2),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba75ab8),
	.w1(32'hbc0e8dba),
	.w2(32'h3c558d09),
	.w3(32'h3bda5f86),
	.w4(32'hbbb8dea1),
	.w5(32'h3b891189),
	.w6(32'hbb044eca),
	.w7(32'h3beae0c8),
	.w8(32'h3be06150),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af2833e),
	.w1(32'hba43e824),
	.w2(32'hbb9a57ff),
	.w3(32'h3c14a973),
	.w4(32'hb8af534e),
	.w5(32'hbc2bb94d),
	.w6(32'h3be9bd9d),
	.w7(32'hbbc4596f),
	.w8(32'hbc139417),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3fc3ee),
	.w1(32'hbba94c7c),
	.w2(32'hbb21f96a),
	.w3(32'hbc509a3c),
	.w4(32'hb9f85876),
	.w5(32'hbb276823),
	.w6(32'hbbac511f),
	.w7(32'hbaf6053a),
	.w8(32'hba33563b),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc3b8ab),
	.w1(32'hba4de59a),
	.w2(32'h3c4522af),
	.w3(32'hbb71e664),
	.w4(32'hbc3fe0a4),
	.w5(32'hbb81a11e),
	.w6(32'hbb9f728a),
	.w7(32'h3b33eeff),
	.w8(32'h3bce5291),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2fa994),
	.w1(32'hbc4c5888),
	.w2(32'hbbe88a5e),
	.w3(32'h399c94d0),
	.w4(32'hbb9d44cf),
	.w5(32'hbb6a478e),
	.w6(32'hbc7a79ee),
	.w7(32'hbc116c0c),
	.w8(32'hbbe772c3),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b836329),
	.w1(32'h3be03141),
	.w2(32'h3b8e1b2e),
	.w3(32'hba6ce7bd),
	.w4(32'h3bff0add),
	.w5(32'h3bcac073),
	.w6(32'h3c3b1827),
	.w7(32'h3c1ba9f8),
	.w8(32'hbb4cb833),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8711e4c),
	.w1(32'h3ac41103),
	.w2(32'hb9c4f01d),
	.w3(32'hbbe0adb3),
	.w4(32'h3a10147b),
	.w5(32'hbab55e34),
	.w6(32'hbb5a1764),
	.w7(32'hb9d9f743),
	.w8(32'hba942dfa),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38feb2b3),
	.w1(32'hbada6ddc),
	.w2(32'hbbbbd3db),
	.w3(32'h3b2946af),
	.w4(32'hbbab5c18),
	.w5(32'hbb4dd06e),
	.w6(32'h3b88f45e),
	.w7(32'hbbc01a5d),
	.w8(32'hbbafef3f),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8e2941),
	.w1(32'hbb29a9f8),
	.w2(32'hbbbc3fc8),
	.w3(32'h3a64e927),
	.w4(32'hbbe4d439),
	.w5(32'hbbf75780),
	.w6(32'h3b5008a8),
	.w7(32'hbb9bdf27),
	.w8(32'hbbe352cb),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb570460),
	.w1(32'hba89157d),
	.w2(32'hbabf12d0),
	.w3(32'hb9cb232a),
	.w4(32'hbaf9d1ab),
	.w5(32'h3ae9362c),
	.w6(32'hb9d8e958),
	.w7(32'hba4273dd),
	.w8(32'hb854bfd4),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b32410),
	.w1(32'hbac3f895),
	.w2(32'h3bde5a6d),
	.w3(32'h3b864489),
	.w4(32'h3b882fca),
	.w5(32'h3cb6c882),
	.w6(32'h3afc37cd),
	.w7(32'h3b30f362),
	.w8(32'h3cc22aa7),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb40e85),
	.w1(32'h3c1139e3),
	.w2(32'hbc231895),
	.w3(32'h3c7f8d99),
	.w4(32'hbbe0984a),
	.w5(32'hbbd87ea2),
	.w6(32'h3bd77c9d),
	.w7(32'hbbe6b9e5),
	.w8(32'hbb89a7ca),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba72bb61),
	.w1(32'hbbe0eda2),
	.w2(32'hbb73600e),
	.w3(32'hbb801b13),
	.w4(32'hbb0e4fc2),
	.w5(32'hbabf0d7a),
	.w6(32'hbbd31cc5),
	.w7(32'hbb83e6b1),
	.w8(32'hbbb66d75),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb46d207),
	.w1(32'hbc03e9cc),
	.w2(32'hbc2f6bf6),
	.w3(32'hbc21844e),
	.w4(32'hbc2308d8),
	.w5(32'hbc751e4a),
	.w6(32'hbc431c92),
	.w7(32'hbba8eb7d),
	.w8(32'hbc6f0c60),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbea68b1),
	.w1(32'hbc81352d),
	.w2(32'h3a6c018d),
	.w3(32'h3b83ab6c),
	.w4(32'h3b80bbe8),
	.w5(32'hbb80c5b8),
	.w6(32'hbb517a2e),
	.w7(32'h3a6d83c6),
	.w8(32'hbaff11cd),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0bc5e5),
	.w1(32'hbbc8835f),
	.w2(32'hbb791ad0),
	.w3(32'hbbef6ad5),
	.w4(32'h3ab68181),
	.w5(32'h3b1f8b84),
	.w6(32'hbb0ad4c6),
	.w7(32'h3a661bcb),
	.w8(32'h3b878bcf),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfda434),
	.w1(32'h39db8398),
	.w2(32'hbc09808c),
	.w3(32'hbb98ed6a),
	.w4(32'hbbb58ae0),
	.w5(32'hbc32729e),
	.w6(32'h3a425475),
	.w7(32'hbbddd213),
	.w8(32'hbc34b60e),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4634e3),
	.w1(32'hbc057ae8),
	.w2(32'hbb87c324),
	.w3(32'hbbcb18fe),
	.w4(32'hbbb90d5f),
	.w5(32'h3b396c9d),
	.w6(32'hbbda289c),
	.w7(32'hbb8aafb0),
	.w8(32'h3b521d38),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa7ada1),
	.w1(32'hbb2bf1ef),
	.w2(32'hbb408e08),
	.w3(32'h3a0ec226),
	.w4(32'hbb6e5e2d),
	.w5(32'hbc0282b4),
	.w6(32'hb86d0650),
	.w7(32'hbb441e05),
	.w8(32'hbbc7c17c),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd69639),
	.w1(32'hbb941137),
	.w2(32'hba8dbde7),
	.w3(32'hbadf1cbc),
	.w4(32'h3ae63c09),
	.w5(32'h3b41ee9d),
	.w6(32'h3a37ba3a),
	.w7(32'h3ac8ab95),
	.w8(32'h3b2f1057),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a44f434),
	.w1(32'h3adfc728),
	.w2(32'hbb89f24f),
	.w3(32'hbb9d8624),
	.w4(32'hbb9f3b18),
	.w5(32'h3b5c5718),
	.w6(32'hbb89c414),
	.w7(32'hbb8a224e),
	.w8(32'h3b206507),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad52ad6),
	.w1(32'hbb105caa),
	.w2(32'hbbcd8371),
	.w3(32'h3c121fe7),
	.w4(32'hbb837ef1),
	.w5(32'hbaf9b56f),
	.w6(32'h3b6418a3),
	.w7(32'hbbcb185d),
	.w8(32'hb926f7d9),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd0f846),
	.w1(32'hbb4fb623),
	.w2(32'hba903d83),
	.w3(32'hbc2f30e4),
	.w4(32'h3ae697c6),
	.w5(32'hbbadf998),
	.w6(32'hbbdc0f41),
	.w7(32'hbb81d651),
	.w8(32'hbc567709),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1c89d5),
	.w1(32'hbba5dbc5),
	.w2(32'hbb806765),
	.w3(32'hbbe45288),
	.w4(32'hbb632e63),
	.w5(32'hbbc14272),
	.w6(32'hbc0d7603),
	.w7(32'hba585e28),
	.w8(32'hbb86fae4),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba5fe71),
	.w1(32'hbaf8f566),
	.w2(32'hbaededf1),
	.w3(32'h3baa6cd4),
	.w4(32'hbae5eea6),
	.w5(32'hba6335f1),
	.w6(32'h3bc3bfbf),
	.w7(32'hbaa3e6d0),
	.w8(32'hba3a1c1c),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b02da16),
	.w1(32'hb9c34a98),
	.w2(32'hb9f6a45b),
	.w3(32'h3b139cc0),
	.w4(32'hbb72bd5e),
	.w5(32'hbbc2c770),
	.w6(32'h3b38d4fb),
	.w7(32'hbbb453e0),
	.w8(32'hbbd86ec5),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1b48d1),
	.w1(32'h3b36e5e2),
	.w2(32'h3b192a7b),
	.w3(32'h3b8be47f),
	.w4(32'h3b1975d3),
	.w5(32'hbc4a70e6),
	.w6(32'h3c1184bf),
	.w7(32'h3b956c3b),
	.w8(32'hbb7b8de7),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b9b63),
	.w1(32'hbbf3a867),
	.w2(32'h3a5d1e52),
	.w3(32'hbbcbad64),
	.w4(32'h3b80b3c1),
	.w5(32'h3c8e0e3e),
	.w6(32'hbc10efe6),
	.w7(32'h3b8970e4),
	.w8(32'h3ca9dd7c),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc01a75),
	.w1(32'h3be9e659),
	.w2(32'h3bbcd21c),
	.w3(32'h3bf879e0),
	.w4(32'h3bf8ea4c),
	.w5(32'h3a939421),
	.w6(32'h3c020f56),
	.w7(32'h3bc4b910),
	.w8(32'h3aa702ca),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0047b0),
	.w1(32'h3b504086),
	.w2(32'h3ad8e5f8),
	.w3(32'h3b1877eb),
	.w4(32'h3b906f85),
	.w5(32'hbc178904),
	.w6(32'h3b561a1a),
	.w7(32'h3bed1e9c),
	.w8(32'hbb60d3c7),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc378ab0),
	.w1(32'hbc0fb88c),
	.w2(32'hbb90cb15),
	.w3(32'hbc0d7a96),
	.w4(32'h3a62586c),
	.w5(32'hbb34e278),
	.w6(32'hbbfe59e6),
	.w7(32'hbb063fc1),
	.w8(32'h3a897426),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba713c1b),
	.w1(32'h3984144f),
	.w2(32'h3a8e0d9d),
	.w3(32'hbb512f92),
	.w4(32'h3acaa52e),
	.w5(32'hbc10466d),
	.w6(32'hbc0f9d92),
	.w7(32'h3a4f91d9),
	.w8(32'hbc0ad397),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1f6fd0),
	.w1(32'hb9a310e4),
	.w2(32'hbb56ee41),
	.w3(32'hbba35630),
	.w4(32'hbb879d44),
	.w5(32'h3b036a4f),
	.w6(32'hbb0e8d5d),
	.w7(32'hbb9c3f3a),
	.w8(32'h3a8d5125),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3812333c),
	.w1(32'hbb79bc95),
	.w2(32'h39a3e059),
	.w3(32'hbc110e92),
	.w4(32'hba01feab),
	.w5(32'hb9e28fa3),
	.w6(32'hbbdf94d0),
	.w7(32'h39d024b9),
	.w8(32'hbb1fa270),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab6f766),
	.w1(32'h3af5dff2),
	.w2(32'hbb939027),
	.w3(32'h3b6703f9),
	.w4(32'hbb953d5d),
	.w5(32'h3b76209e),
	.w6(32'h3b7bce87),
	.w7(32'hbbf0612d),
	.w8(32'h3b994c01),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397ba69e),
	.w1(32'hbbe6bde7),
	.w2(32'hbb66fa77),
	.w3(32'h3bc9979e),
	.w4(32'hbb73a191),
	.w5(32'hbc125a17),
	.w6(32'hbbab11c2),
	.w7(32'hbbb3f56c),
	.w8(32'hbc601be2),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb88248b),
	.w1(32'hbc0cc734),
	.w2(32'hba8777c4),
	.w3(32'hbc11d3c2),
	.w4(32'h3b7f2387),
	.w5(32'hbaf77948),
	.w6(32'hbc34a1c4),
	.w7(32'hbb92315f),
	.w8(32'hbb433bfa),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0afe21),
	.w1(32'h3b4ed069),
	.w2(32'hb91133ac),
	.w3(32'hbb9e04bc),
	.w4(32'h39b1c070),
	.w5(32'hbb0ed244),
	.w6(32'hbb95e63b),
	.w7(32'hb9a326b8),
	.w8(32'hbac1f23c),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb06375e),
	.w1(32'h3a840479),
	.w2(32'hbb05669f),
	.w3(32'hb8ff3432),
	.w4(32'hb99339b0),
	.w5(32'hb9e298a9),
	.w6(32'h38206eb6),
	.w7(32'hbb1ef6c4),
	.w8(32'h3b61d813),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7166c9),
	.w1(32'h3bbde903),
	.w2(32'h3ae9c3a1),
	.w3(32'hbb80fddf),
	.w4(32'hbb0d0a2f),
	.w5(32'hbb46719e),
	.w6(32'h39844c7b),
	.w7(32'hbaeefec7),
	.w8(32'hbbdcf2d1),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb448e40),
	.w1(32'hbbd630b4),
	.w2(32'hbb134e35),
	.w3(32'hbc29eb07),
	.w4(32'h3b0165ee),
	.w5(32'hbbb6cb74),
	.w6(32'hbc29516c),
	.w7(32'h3af6f1a7),
	.w8(32'hbc30443f),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc061e3f),
	.w1(32'hbbe4f2ba),
	.w2(32'hbb4d600a),
	.w3(32'hbb94de0d),
	.w4(32'h3a0491f5),
	.w5(32'hbbe2d594),
	.w6(32'hbc077edd),
	.w7(32'hbc03e812),
	.w8(32'hbc2d6553),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb985a8f),
	.w1(32'h3b1ec03b),
	.w2(32'h3abb12a8),
	.w3(32'hbb80faa3),
	.w4(32'h3b479cb1),
	.w5(32'h3b877132),
	.w6(32'hbbc98485),
	.w7(32'h3b5cc258),
	.w8(32'h3b84a245),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8d7058),
	.w1(32'hbbcaa082),
	.w2(32'hbbca50fe),
	.w3(32'h3b3976ca),
	.w4(32'hbbe9a146),
	.w5(32'h3bd03106),
	.w6(32'hba229fc9),
	.w7(32'hbbfd2d32),
	.w8(32'h3b91b9f2),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8c6a64),
	.w1(32'h3c020b66),
	.w2(32'h3bd4066c),
	.w3(32'h3c6ea990),
	.w4(32'h3bb70528),
	.w5(32'h39d5d106),
	.w6(32'h3c5c3785),
	.w7(32'hbae365b5),
	.w8(32'hbbd84638),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba621b01),
	.w1(32'hbbc6389b),
	.w2(32'h3ca8651d),
	.w3(32'hba643896),
	.w4(32'h3c8f0f7d),
	.w5(32'h3d02d062),
	.w6(32'hbc0eb288),
	.w7(32'h3ca72453),
	.w8(32'h3cf66065),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd3f803),
	.w1(32'h3bdca533),
	.w2(32'hba38b211),
	.w3(32'h3c0f003b),
	.w4(32'hbaa5001d),
	.w5(32'h3a39e28a),
	.w6(32'h3b7d7f06),
	.w7(32'hbb5eb608),
	.w8(32'hbab91a59),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacd9a7a),
	.w1(32'h3b40a30d),
	.w2(32'hbb099485),
	.w3(32'h3b077237),
	.w4(32'hb99bd957),
	.w5(32'hbb192574),
	.w6(32'h3bca88b5),
	.w7(32'hbaae230c),
	.w8(32'hbb2b19a4),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1f1125),
	.w1(32'h3ad4ee36),
	.w2(32'hba981660),
	.w3(32'h3ac31cc1),
	.w4(32'h3ad1e7c3),
	.w5(32'hbbb06289),
	.w6(32'h3b415876),
	.w7(32'h39e8b9dd),
	.w8(32'hbaf1c680),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb61faba),
	.w1(32'h3bb245ad),
	.w2(32'hbbb5f5da),
	.w3(32'h3ad33595),
	.w4(32'hbb83c8c3),
	.w5(32'hba8d642a),
	.w6(32'hba6990bc),
	.w7(32'hbbce678d),
	.w8(32'hbb30b66f),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2c92ac),
	.w1(32'hbbbfd414),
	.w2(32'h3b14c5c8),
	.w3(32'hbbbfd0e8),
	.w4(32'hbb28af81),
	.w5(32'h3b0d3165),
	.w6(32'hbbfb6ec3),
	.w7(32'h3aad006c),
	.w8(32'h3c13d83c),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba97250e),
	.w1(32'hbb8e7657),
	.w2(32'hbbf445d2),
	.w3(32'h3bc7ccc5),
	.w4(32'hb9c869fb),
	.w5(32'hbbc5b207),
	.w6(32'h3b826420),
	.w7(32'hbb44b79b),
	.w8(32'hbc011284),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc48efdf),
	.w1(32'hbba2225d),
	.w2(32'hba506f2d),
	.w3(32'hbbf1b14a),
	.w4(32'hba2a601c),
	.w5(32'hbaa2bc99),
	.w6(32'hbbe445c4),
	.w7(32'hba4837f2),
	.w8(32'hb935dfec),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba914f3b),
	.w1(32'h3afca56d),
	.w2(32'hbbd09328),
	.w3(32'h3aabcd5e),
	.w4(32'hbb5fed9e),
	.w5(32'hbb73e441),
	.w6(32'h3b13599e),
	.w7(32'hbbebdc21),
	.w8(32'hbc0cdcb0),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc192e35),
	.w1(32'hbba32319),
	.w2(32'h3bc214b6),
	.w3(32'hbbf0343d),
	.w4(32'hb9bd5ce1),
	.w5(32'h390ac457),
	.w6(32'hbbf27853),
	.w7(32'h3bdc3bae),
	.w8(32'h3a9a3975),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36f56d29),
	.w1(32'hbc0ba4dd),
	.w2(32'hbaeaf7e3),
	.w3(32'hbc6b42d0),
	.w4(32'h3a1bd999),
	.w5(32'h3c03190f),
	.w6(32'hbc9fd64f),
	.w7(32'hbb03fb1e),
	.w8(32'h3c07787f),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b87496f),
	.w1(32'h3c05fe29),
	.w2(32'hbc135da8),
	.w3(32'h3b915392),
	.w4(32'hbb94c1de),
	.w5(32'h3b541a55),
	.w6(32'h3c127dfd),
	.w7(32'hbba1385b),
	.w8(32'h3ad34826),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9fce22),
	.w1(32'h3ba5adc0),
	.w2(32'hbb4586e8),
	.w3(32'h3a355864),
	.w4(32'hbaadbb4d),
	.w5(32'hbb786a80),
	.w6(32'h3938a33a),
	.w7(32'hbb3f513b),
	.w8(32'hbb0d4b43),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule