module layer_8_featuremap_31(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d0899c),
	.w1(32'hba22c394),
	.w2(32'hb8a0560b),
	.w3(32'hba82b27c),
	.w4(32'hb8124427),
	.w5(32'hb89317f6),
	.w6(32'hb8efaec3),
	.w7(32'hb9736887),
	.w8(32'hb9bc7157),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e9a868),
	.w1(32'hb9ea10ed),
	.w2(32'hb9901db8),
	.w3(32'hba2e942e),
	.w4(32'hb9c55f7e),
	.w5(32'hb98d957a),
	.w6(32'hb99a6f7f),
	.w7(32'hb9cefe68),
	.w8(32'h39c2025f),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb81b932b),
	.w1(32'hb97d7938),
	.w2(32'hb8b45bd7),
	.w3(32'hb95d2838),
	.w4(32'h3789d087),
	.w5(32'h3960a138),
	.w6(32'h38f1fe9c),
	.w7(32'hb897bdb8),
	.w8(32'hbab38fb9),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f3edb4),
	.w1(32'hbb095936),
	.w2(32'hb9ce0c43),
	.w3(32'h3a5cbfbf),
	.w4(32'hbaec2b77),
	.w5(32'hbaad8e6d),
	.w6(32'hb9034ab5),
	.w7(32'h39838f96),
	.w8(32'h392e7b69),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fbb109),
	.w1(32'hb988c2ce),
	.w2(32'hb8b50a4b),
	.w3(32'hba1fdbc7),
	.w4(32'h38306ab7),
	.w5(32'h37b32e65),
	.w6(32'h3974d8ea),
	.w7(32'h3971a67b),
	.w8(32'h3a89b825),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae87498),
	.w1(32'h39e49fa0),
	.w2(32'h3b0cbcfa),
	.w3(32'h3aba71e5),
	.w4(32'h3a3ada05),
	.w5(32'h3aae6af0),
	.w6(32'h3ab0c2b8),
	.w7(32'h3b3b6e2a),
	.w8(32'h3a2fb522),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9980ebd),
	.w1(32'hb9e4a967),
	.w2(32'hb9ae2a8b),
	.w3(32'hba5237a6),
	.w4(32'hb98b50fd),
	.w5(32'h3898fc51),
	.w6(32'h373ba905),
	.w7(32'hba1be29c),
	.w8(32'hb80ad654),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2cded4),
	.w1(32'hb94f4f90),
	.w2(32'hb868767d),
	.w3(32'hba25657f),
	.w4(32'h383ad772),
	.w5(32'hb94c7e46),
	.w6(32'h39ab454e),
	.w7(32'h39e70b39),
	.w8(32'h39fe0fff),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b13f95),
	.w1(32'hb847962f),
	.w2(32'hb9b2ab9f),
	.w3(32'hba850b4d),
	.w4(32'hb92a3918),
	.w5(32'h390ebb46),
	.w6(32'h3997b0ac),
	.w7(32'hba53d647),
	.w8(32'hbb973efa),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf62282),
	.w1(32'hbab27882),
	.w2(32'hbb7ecfe1),
	.w3(32'hbaaaa707),
	.w4(32'hbb84687c),
	.w5(32'hbaf19321),
	.w6(32'hbbc1e563),
	.w7(32'hb9691b0e),
	.w8(32'h3a24282b),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ab21f8),
	.w1(32'h3927ea6a),
	.w2(32'hb98bbf50),
	.w3(32'hb8d9be25),
	.w4(32'h3a1a5c55),
	.w5(32'h3a109203),
	.w6(32'h3a2da90b),
	.w7(32'h397c9e0c),
	.w8(32'h39bfb248),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9958a07),
	.w1(32'hb9d1deb2),
	.w2(32'h387944b8),
	.w3(32'hba22d31f),
	.w4(32'hb8eb38ac),
	.w5(32'h393ccc0c),
	.w6(32'h392060b2),
	.w7(32'hb7bedb66),
	.w8(32'h3a1f3a3e),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392d3357),
	.w1(32'hb902be72),
	.w2(32'hb9754296),
	.w3(32'h3827b237),
	.w4(32'h38a0d058),
	.w5(32'h390bb795),
	.w6(32'h3a236b5d),
	.w7(32'hb93daff8),
	.w8(32'h3ace02a5),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b06945d),
	.w1(32'h39c3d892),
	.w2(32'h3b1b9f74),
	.w3(32'h3ae3f0cd),
	.w4(32'h3a5df4cb),
	.w5(32'h3acc8122),
	.w6(32'h3ac73c5c),
	.w7(32'h3b515663),
	.w8(32'h3a9eb2aa),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a80177d),
	.w1(32'h39f4b512),
	.w2(32'h3ab39ffb),
	.w3(32'h3a70d518),
	.w4(32'h3a25a16e),
	.w5(32'h3a8f235b),
	.w6(32'h3a77a372),
	.w7(32'h3b07d864),
	.w8(32'hb9c5f953),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99b6d22),
	.w1(32'hb9a52fed),
	.w2(32'hba5d4a64),
	.w3(32'hba179003),
	.w4(32'hb9ec56f5),
	.w5(32'hba25c017),
	.w6(32'hba34b2b9),
	.w7(32'hb9d5123b),
	.w8(32'hbb6ddedf),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad07255),
	.w1(32'hbb583e81),
	.w2(32'hba0473c6),
	.w3(32'hb9e8683a),
	.w4(32'hbab57843),
	.w5(32'hbb01a4fa),
	.w6(32'hbb3ded5c),
	.w7(32'hbafe999d),
	.w8(32'h3912bf86),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb961626e),
	.w1(32'hba740749),
	.w2(32'hba42107b),
	.w3(32'hba3b6d2a),
	.w4(32'hb92c7de1),
	.w5(32'hba0d747b),
	.w6(32'h3950e53a),
	.w7(32'hba15441c),
	.w8(32'hba3e7066),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba459846),
	.w1(32'h3a2bcfd6),
	.w2(32'h3a3957dc),
	.w3(32'hb9e2b794),
	.w4(32'h3a73044c),
	.w5(32'h395fd1c6),
	.w6(32'h3ac7f505),
	.w7(32'h3ab80389),
	.w8(32'hbbae056f),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2fb16c),
	.w1(32'hbbb00107),
	.w2(32'hbb183f22),
	.w3(32'hbb4967d5),
	.w4(32'hbb8722c6),
	.w5(32'hbb432824),
	.w6(32'hbbc6d6cb),
	.w7(32'hbbaed1c1),
	.w8(32'h3a95939b),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a68abf5),
	.w1(32'h3a67a5b3),
	.w2(32'h3a0f822e),
	.w3(32'h3a99b6fe),
	.w4(32'h3a912bd9),
	.w5(32'h3ad1cdc4),
	.w6(32'h3a3e0654),
	.w7(32'hb883ea69),
	.w8(32'h3a1eca88),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba39c4a3),
	.w1(32'hba3d4667),
	.w2(32'h39a5b59d),
	.w3(32'hba8a3b0e),
	.w4(32'hb953a364),
	.w5(32'h3a5d56f9),
	.w6(32'h3999aa4d),
	.w7(32'h39c424bc),
	.w8(32'h3acedb6e),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3934463b),
	.w1(32'hba30f7fb),
	.w2(32'hba94a7ae),
	.w3(32'h3a643a18),
	.w4(32'h387abf2c),
	.w5(32'hb93e0a59),
	.w6(32'hba1e313e),
	.w7(32'hbb03e5d4),
	.w8(32'hb9caa04b),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96786a6),
	.w1(32'hb7d6e00e),
	.w2(32'h38f6eb9a),
	.w3(32'hb99eb75c),
	.w4(32'h3a01da86),
	.w5(32'hba82d633),
	.w6(32'h3a79e5b0),
	.w7(32'h39d60092),
	.w8(32'hbb3b73ad),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0ba579),
	.w1(32'hba4f8f1a),
	.w2(32'hbab39b98),
	.w3(32'hbb291c2f),
	.w4(32'hbb1c96d4),
	.w5(32'hbb0fddd1),
	.w6(32'hbb06c5d5),
	.w7(32'hbb0b9ad1),
	.w8(32'h3a92ea19),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390026c4),
	.w1(32'hb9d6a65f),
	.w2(32'hba5443b7),
	.w3(32'h3a744db4),
	.w4(32'h39981b96),
	.w5(32'h392f92fb),
	.w6(32'hb984c574),
	.w7(32'hbac93cdd),
	.w8(32'h3a531433),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f3ecbf),
	.w1(32'hb9ae3921),
	.w2(32'hba3faa50),
	.w3(32'h3a49d00d),
	.w4(32'h395e415c),
	.w5(32'h38bc8220),
	.w6(32'hb99226e4),
	.w7(32'hbab1317b),
	.w8(32'h39aa8069),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f5f44c),
	.w1(32'hb9faefab),
	.w2(32'hb8b0d878),
	.w3(32'hb92965be),
	.w4(32'h382e280d),
	.w5(32'h39b6afc2),
	.w6(32'h39a357d0),
	.w7(32'hba4e6e8d),
	.w8(32'hbb29ec56),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba368e3a),
	.w1(32'h3aa172b3),
	.w2(32'hbb4103a3),
	.w3(32'hbabfcb59),
	.w4(32'hb925ff8a),
	.w5(32'hbb3eeef1),
	.w6(32'hbbae7153),
	.w7(32'hb9d5a9be),
	.w8(32'h395a6f5d),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91fb354),
	.w1(32'hb9533cb1),
	.w2(32'hb75515af),
	.w3(32'hb975c745),
	.w4(32'hb7a0c37b),
	.w5(32'h38e9f2fa),
	.w6(32'h39104187),
	.w7(32'h395d48a3),
	.w8(32'hbaaa3d36),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab564dd),
	.w1(32'hba605d40),
	.w2(32'h3b75615f),
	.w3(32'h3a3bb73e),
	.w4(32'h3a21e5fc),
	.w5(32'hb9f8caec),
	.w6(32'hbb20dc66),
	.w7(32'hba6825e8),
	.w8(32'h3adf49c7),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99ecbcd),
	.w1(32'h3a24317d),
	.w2(32'hba4e2497),
	.w3(32'hb86b1bc2),
	.w4(32'h3ae29823),
	.w5(32'h3af92876),
	.w6(32'h39b4777e),
	.w7(32'hbae553cf),
	.w8(32'hba7d27c0),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb02577b),
	.w1(32'hbbaea63c),
	.w2(32'hbb144da3),
	.w3(32'hbafea506),
	.w4(32'hbb512770),
	.w5(32'hbb880576),
	.w6(32'hbad01abf),
	.w7(32'h3a0585c8),
	.w8(32'h3affa1f1),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8d00a3),
	.w1(32'h3b062df6),
	.w2(32'h3ae15e86),
	.w3(32'h3aa6b3cb),
	.w4(32'hba9f12ed),
	.w5(32'h39f21499),
	.w6(32'h3bc1029f),
	.w7(32'h3b6f5e15),
	.w8(32'h3aa6e522),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad910e8),
	.w1(32'h3965a9ba),
	.w2(32'h3b01a43a),
	.w3(32'h3ab4bb83),
	.w4(32'h3a27aa54),
	.w5(32'h3aa3f543),
	.w6(32'h3aa1a200),
	.w7(32'h3b35df7e),
	.w8(32'hb95a7ec3),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cb3791),
	.w1(32'h388ecbca),
	.w2(32'h39a73f1b),
	.w3(32'hba274cce),
	.w4(32'h39deda28),
	.w5(32'hb9f06d1c),
	.w6(32'h3a424668),
	.w7(32'h399ed643),
	.w8(32'h3a125b79),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba52dfc6),
	.w1(32'hba387e8f),
	.w2(32'hba458452),
	.w3(32'hb9cd101d),
	.w4(32'hba892508),
	.w5(32'hb9f3cb6c),
	.w6(32'h38b3fa4a),
	.w7(32'hba81358a),
	.w8(32'h39fc3fad),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h373a14b4),
	.w1(32'hb980e9dd),
	.w2(32'h39ab7eaf),
	.w3(32'hb8c4e9c0),
	.w4(32'h398862a5),
	.w5(32'h3a1e5f06),
	.w6(32'h39c54d77),
	.w7(32'h3a05798b),
	.w8(32'h3b1caa56),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b01bab9),
	.w1(32'h3a8681b7),
	.w2(32'h3b2cc867),
	.w3(32'h3b1dad5d),
	.w4(32'h3aaf9d60),
	.w5(32'h3b0b3aad),
	.w6(32'h3b034e2f),
	.w7(32'h3b88f0ec),
	.w8(32'h38457597),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2fabb6),
	.w1(32'hba5590cb),
	.w2(32'hba81a397),
	.w3(32'hba251563),
	.w4(32'hba21a3b3),
	.w5(32'hb9c4f097),
	.w6(32'hba94ae6a),
	.w7(32'hbabda7d5),
	.w8(32'h3987422b),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7651ac6),
	.w1(32'hb9841b94),
	.w2(32'hb9e2f911),
	.w3(32'h39cb87b8),
	.w4(32'h3902b783),
	.w5(32'h37e1c191),
	.w6(32'hb8d3ee17),
	.w7(32'hba2a87f6),
	.w8(32'h3bac1d36),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2932e6),
	.w1(32'hbb7113cc),
	.w2(32'hbbbc6e16),
	.w3(32'h3b2bb5c1),
	.w4(32'h3bb61d16),
	.w5(32'h3a6f86b1),
	.w6(32'hba86b746),
	.w7(32'hbaaeb1bc),
	.w8(32'hbc37a224),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaca1096),
	.w1(32'hbc448859),
	.w2(32'h3cda1f84),
	.w3(32'hbc0c1ce5),
	.w4(32'hbc0566bc),
	.w5(32'h3bd82a8b),
	.w6(32'h3afa9ac3),
	.w7(32'h37beaec9),
	.w8(32'h3b414a95),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7536cd),
	.w1(32'hbbab3ea0),
	.w2(32'hbb7ed6f1),
	.w3(32'h3b1822b4),
	.w4(32'hba32279a),
	.w5(32'hbafb95fd),
	.w6(32'hbb05950b),
	.w7(32'hbba0127e),
	.w8(32'h3b71ce8c),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2483ac),
	.w1(32'hbb892bf6),
	.w2(32'hbb8dbf30),
	.w3(32'h3b8ec94f),
	.w4(32'h3a3ce611),
	.w5(32'hbbc84f86),
	.w6(32'hba983ffe),
	.w7(32'hbb4f68b8),
	.w8(32'hbb0bae9d),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb37c8e9),
	.w1(32'h3b699416),
	.w2(32'hbba33ff8),
	.w3(32'hbbf7dc47),
	.w4(32'hbbb0d3dc),
	.w5(32'hbabc3523),
	.w6(32'hbc003178),
	.w7(32'hbb7d0079),
	.w8(32'hbbf860ae),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc829342),
	.w1(32'h3d115cc1),
	.w2(32'hbb024817),
	.w3(32'hbb8a0637),
	.w4(32'hbcab8fd9),
	.w5(32'hba989060),
	.w6(32'h3c60ec21),
	.w7(32'h3c4514a9),
	.w8(32'hbbc851bf),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388ebead),
	.w1(32'hbb95a3a2),
	.w2(32'h3a3f73bc),
	.w3(32'h3ba64463),
	.w4(32'h3b3789e2),
	.w5(32'h3b974d43),
	.w6(32'hbbc4afe1),
	.w7(32'h3bb9ddbf),
	.w8(32'h39300d60),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdf4a10),
	.w1(32'h3b08a387),
	.w2(32'h3c202087),
	.w3(32'hbbadb921),
	.w4(32'h3b3394ac),
	.w5(32'h3c3b9954),
	.w6(32'h3bbe6097),
	.w7(32'h3c89e873),
	.w8(32'h3af5e3de),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aac7c39),
	.w1(32'hbc11b76d),
	.w2(32'hbb84713a),
	.w3(32'h3b2e06c7),
	.w4(32'hba37bf63),
	.w5(32'hbb0b8a73),
	.w6(32'hbbb9f10a),
	.w7(32'hba5f9133),
	.w8(32'h3a838460),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acd1567),
	.w1(32'hbb550926),
	.w2(32'hbb8218e6),
	.w3(32'h3b1b917b),
	.w4(32'hbb286704),
	.w5(32'hbba21f63),
	.w6(32'hbb476f02),
	.w7(32'hbbc23e5f),
	.w8(32'h3bc07faf),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdbebee),
	.w1(32'hbbed2f86),
	.w2(32'hbc07ba62),
	.w3(32'h3bc176a6),
	.w4(32'hbb5f6306),
	.w5(32'hbc1c1f77),
	.w6(32'hbbc48bdf),
	.w7(32'hbc51ef87),
	.w8(32'h3c9f804c),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c906e5b),
	.w1(32'hbb3dc3d5),
	.w2(32'h3bac1fb0),
	.w3(32'h3c98608b),
	.w4(32'hbbb69a68),
	.w5(32'h3b47fa8c),
	.w6(32'hbb5f1aa6),
	.w7(32'hbb0985b8),
	.w8(32'hbb9c0192),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb997b1a),
	.w1(32'hba96f38d),
	.w2(32'h388c4afc),
	.w3(32'hbb44e201),
	.w4(32'hb895c106),
	.w5(32'hbb276234),
	.w6(32'h3ac1f96e),
	.w7(32'h3c1801dc),
	.w8(32'h3c01f872),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd40681),
	.w1(32'h3cf5170b),
	.w2(32'hbbab6276),
	.w3(32'h3c2ac1f2),
	.w4(32'h3cc1bda0),
	.w5(32'hbc766223),
	.w6(32'h3d16a66a),
	.w7(32'h3b07c8c9),
	.w8(32'hbbd8c950),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9dc81f),
	.w1(32'hbc022b9f),
	.w2(32'hbc8e90fa),
	.w3(32'hbc277770),
	.w4(32'h3ae4a3ae),
	.w5(32'hbbccad32),
	.w6(32'hbb375c42),
	.w7(32'hbc080dbb),
	.w8(32'hbc48c217),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb310efb),
	.w1(32'hbb0c2a74),
	.w2(32'h3b2586d8),
	.w3(32'hbba72c3c),
	.w4(32'hbc20b64d),
	.w5(32'h3bb10a80),
	.w6(32'hbba00e34),
	.w7(32'hba962a9a),
	.w8(32'h3bd22b2f),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc70373d),
	.w1(32'h3d5300b5),
	.w2(32'hbb0a9801),
	.w3(32'hbc8544e6),
	.w4(32'h3c1076b8),
	.w5(32'h3c8e0fa1),
	.w6(32'hbac02a84),
	.w7(32'hbc8be572),
	.w8(32'h3c41c631),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf044d3),
	.w1(32'hbb93bb2c),
	.w2(32'h3ad8fb51),
	.w3(32'h3c261d11),
	.w4(32'h39ffbeb7),
	.w5(32'h3b304773),
	.w6(32'h3ae551ae),
	.w7(32'h3b8bf655),
	.w8(32'h3b888409),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b84ce33),
	.w1(32'h3b88452e),
	.w2(32'h3a3a3356),
	.w3(32'h3b48efb0),
	.w4(32'h3bfa4427),
	.w5(32'hbbd310f5),
	.w6(32'h39def511),
	.w7(32'hba36fd4a),
	.w8(32'hbc85116f),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbceed0e7),
	.w1(32'h3c4517e4),
	.w2(32'h3c0b6f80),
	.w3(32'hbc88ce0c),
	.w4(32'hbbb6036e),
	.w5(32'hbbd31ea6),
	.w6(32'hbd04030a),
	.w7(32'hbc0f9a27),
	.w8(32'hbb1ee53a),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb763438),
	.w1(32'h3a9022c1),
	.w2(32'hbbd1d610),
	.w3(32'h3b037e82),
	.w4(32'hbb8ab675),
	.w5(32'hbb0349dc),
	.w6(32'hbb4d0b5c),
	.w7(32'hb9a6bd4d),
	.w8(32'h3b30760f),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a72f35a),
	.w1(32'hbc85ea20),
	.w2(32'hbc3107f8),
	.w3(32'h3a6a6b40),
	.w4(32'hbc36f130),
	.w5(32'hbc69ebf3),
	.w6(32'hbc257c25),
	.w7(32'hbc279f09),
	.w8(32'hb73b7cd5),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1b2216),
	.w1(32'h3cc58bf7),
	.w2(32'h3d00e4ba),
	.w3(32'hbc0a0296),
	.w4(32'hbca90c2e),
	.w5(32'h3a0e47a3),
	.w6(32'h3c4cd94b),
	.w7(32'hb9364c9f),
	.w8(32'h3afa86d1),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8f4b83),
	.w1(32'hbb281dfb),
	.w2(32'hba0fee1a),
	.w3(32'h3aa3a6f5),
	.w4(32'hb9e26cec),
	.w5(32'hbab2383a),
	.w6(32'hba1d3840),
	.w7(32'hbae30e7f),
	.w8(32'h3b5e27d2),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7b6648),
	.w1(32'hbac5b005),
	.w2(32'hba085bdc),
	.w3(32'h3b5a51cd),
	.w4(32'h3a8ad1c5),
	.w5(32'hba91682a),
	.w6(32'hb9e0ea3d),
	.w7(32'hbb1f88de),
	.w8(32'h3b2f3527),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b384291),
	.w1(32'hbb0e2935),
	.w2(32'hbb316f91),
	.w3(32'h3b227fad),
	.w4(32'hb986e468),
	.w5(32'hbb48a67e),
	.w6(32'hbad42c11),
	.w7(32'hbb95349f),
	.w8(32'h3ac7fecc),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc267765),
	.w1(32'h3b416aac),
	.w2(32'hbc20a371),
	.w3(32'hbb24a476),
	.w4(32'hbb7f61fb),
	.w5(32'hba054935),
	.w6(32'h3b505de0),
	.w7(32'hbbe6fad5),
	.w8(32'h3a9dcc1d),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b94f78),
	.w1(32'hbbbdc06c),
	.w2(32'hbb917efa),
	.w3(32'h3ab47c0d),
	.w4(32'hbace546a),
	.w5(32'hbb39775e),
	.w6(32'hbb820b9c),
	.w7(32'hbb0b660e),
	.w8(32'h3c9eb90a),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca45529),
	.w1(32'hbc0a3618),
	.w2(32'hbc101b0e),
	.w3(32'h3cb8738c),
	.w4(32'hbb22c9e6),
	.w5(32'hbc12be6e),
	.w6(32'hbb0e10d5),
	.w7(32'hbc38a03a),
	.w8(32'h3c0dd25c),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2ee891),
	.w1(32'hbadbdef0),
	.w2(32'hbb470155),
	.w3(32'h3bd986bf),
	.w4(32'h3b887b52),
	.w5(32'hba833c98),
	.w6(32'hb9cc7d77),
	.w7(32'hbb2fb919),
	.w8(32'h39d3795b),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacc73c6),
	.w1(32'hbbe020e2),
	.w2(32'hbb9448ea),
	.w3(32'h39ba36d1),
	.w4(32'hb9c9e452),
	.w5(32'hbabac6d9),
	.w6(32'hbbd600ef),
	.w7(32'hba72628d),
	.w8(32'h3c3e7b7b),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7605d7),
	.w1(32'hbaae27c8),
	.w2(32'hbb81cc87),
	.w3(32'h3c35f7c3),
	.w4(32'h3b9940c8),
	.w5(32'hba45a3d5),
	.w6(32'h377eb1db),
	.w7(32'hbb842553),
	.w8(32'hbc0af439),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c92ae5f),
	.w1(32'hbb8c7764),
	.w2(32'hbc2feb79),
	.w3(32'h3c743214),
	.w4(32'h3c45bcbe),
	.w5(32'hbbe00ba0),
	.w6(32'hbaa7627e),
	.w7(32'hb93720a9),
	.w8(32'h3b7965bf),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e1ebc2),
	.w1(32'h3b1d41c9),
	.w2(32'hbc05d0d3),
	.w3(32'hbb027592),
	.w4(32'h3b10c0cc),
	.w5(32'hbb9da60b),
	.w6(32'hbac9e3ab),
	.w7(32'hbbfacc8c),
	.w8(32'h3bbd472d),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be189da),
	.w1(32'hbb7e0085),
	.w2(32'hbb57a71d),
	.w3(32'h3b8af43b),
	.w4(32'h3ad4dfb1),
	.w5(32'hbb0906c9),
	.w6(32'hbb071865),
	.w7(32'hbb9a4a7e),
	.w8(32'h3bd4cab5),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcc45c3),
	.w1(32'hba8243e6),
	.w2(32'hbba58cec),
	.w3(32'h3ac3d580),
	.w4(32'h3a821cf2),
	.w5(32'hbad30196),
	.w6(32'hba178cdb),
	.w7(32'hbb9ca752),
	.w8(32'h3cc3405b),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc0c3f0),
	.w1(32'hbc21934a),
	.w2(32'hbc1560a6),
	.w3(32'h3cdae438),
	.w4(32'hbb1f3963),
	.w5(32'hbc129654),
	.w6(32'hbad5b79c),
	.w7(32'hbc34f176),
	.w8(32'h3c4039bf),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c89dfe0),
	.w1(32'hbbc22d4a),
	.w2(32'hbbdb7e38),
	.w3(32'h3c88bf83),
	.w4(32'hbb2c8e3a),
	.w5(32'hbb839381),
	.w6(32'hbae870f5),
	.w7(32'hbbb38132),
	.w8(32'hbb21abd7),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcf51e4),
	.w1(32'hba515bca),
	.w2(32'h3b264ee3),
	.w3(32'hbb8200ae),
	.w4(32'hb8886906),
	.w5(32'h3aa767be),
	.w6(32'hbb05d70d),
	.w7(32'h3a9160c7),
	.w8(32'hbcb971ed),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce986e1),
	.w1(32'h38d6b120),
	.w2(32'hbbecd9a6),
	.w3(32'hbb418644),
	.w4(32'hba8add62),
	.w5(32'hbc457b85),
	.w6(32'h3986a1f3),
	.w7(32'hbc0daca4),
	.w8(32'h3ac464e5),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7acc62),
	.w1(32'h3a15305b),
	.w2(32'hbb0092fb),
	.w3(32'h3a14f6a7),
	.w4(32'h39446231),
	.w5(32'hbb633f7c),
	.w6(32'h39f017c0),
	.w7(32'hbbc35514),
	.w8(32'hbc14ccad),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc229722),
	.w1(32'hbb25ebb3),
	.w2(32'hbb0d299c),
	.w3(32'hbbc87d0b),
	.w4(32'hbb9b791a),
	.w5(32'hbb9aaffd),
	.w6(32'hbaf2ef7a),
	.w7(32'hbb2a5f45),
	.w8(32'h3c0777cd),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad7b03b),
	.w1(32'hbbbd6175),
	.w2(32'h3cb5b45d),
	.w3(32'hbb569f31),
	.w4(32'h3c840113),
	.w5(32'hbb12e049),
	.w6(32'hbb943ec3),
	.w7(32'hbc501ecd),
	.w8(32'h3a56daa1),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b228afc),
	.w1(32'hbb8b64e9),
	.w2(32'h3b5b37bb),
	.w3(32'h3b47fcd8),
	.w4(32'hb9a6283d),
	.w5(32'h3bcca293),
	.w6(32'hbb06b6a7),
	.w7(32'h3c00adea),
	.w8(32'h3b087fe6),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a54c384),
	.w1(32'hbc044188),
	.w2(32'hbbd09a1d),
	.w3(32'h3af87b58),
	.w4(32'hbb13c8e7),
	.w5(32'hbbdee5c2),
	.w6(32'hbbc176cb),
	.w7(32'hbba0f966),
	.w8(32'h383b45b5),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc12b89c),
	.w1(32'h3b31f4d9),
	.w2(32'h3c53608a),
	.w3(32'hbbe26499),
	.w4(32'h3b6f6e45),
	.w5(32'h3c78ae20),
	.w6(32'h3bfe0a67),
	.w7(32'h3cb70df2),
	.w8(32'h3b0011b6),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2237d1),
	.w1(32'hbc10ebcd),
	.w2(32'hbac541d7),
	.w3(32'h3ba4b446),
	.w4(32'h3aad9199),
	.w5(32'hb9916c34),
	.w6(32'h3aae6a63),
	.w7(32'hb986693d),
	.w8(32'hbb9dcbe4),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf194b4),
	.w1(32'hbcaba110),
	.w2(32'h3bdaac13),
	.w3(32'hbc04691d),
	.w4(32'hbbc06c80),
	.w5(32'h396b9425),
	.w6(32'hbc5c8d83),
	.w7(32'hbae9d94f),
	.w8(32'h381f3aeb),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0a09cc),
	.w1(32'h3b29f9df),
	.w2(32'h3c463199),
	.w3(32'hbbd537db),
	.w4(32'h3b62a2da),
	.w5(32'h3c696c7d),
	.w6(32'h3beda714),
	.w7(32'h3cab6f8a),
	.w8(32'h38d31499),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe9ed04),
	.w1(32'h3b1686aa),
	.w2(32'h3c2aa132),
	.w3(32'hbbb4e8f2),
	.w4(32'h3b43e11c),
	.w5(32'h3c48a244),
	.w6(32'h3bcef5d1),
	.w7(32'h3c934f23),
	.w8(32'hbba61558),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbccc48c),
	.w1(32'hbbb51696),
	.w2(32'h3ba74327),
	.w3(32'hbb843fcb),
	.w4(32'hbb9886c3),
	.w5(32'h3b0a336c),
	.w6(32'hbb7e223e),
	.w7(32'h3c4adf5d),
	.w8(32'h3b874533),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb328fb4),
	.w1(32'hbb9db05c),
	.w2(32'h3c80576a),
	.w3(32'hbc228b15),
	.w4(32'h3bea928e),
	.w5(32'h3bdf8885),
	.w6(32'hbaa722d5),
	.w7(32'h3c306825),
	.w8(32'h3a877ba7),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399c8ac7),
	.w1(32'hbb1f1de3),
	.w2(32'hbb53d6d9),
	.w3(32'h3a4b345d),
	.w4(32'hbac8d53d),
	.w5(32'hbb669a81),
	.w6(32'hbb24c1aa),
	.w7(32'hbb96d66a),
	.w8(32'h3b8a85a0),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1eb72e),
	.w1(32'h3c872289),
	.w2(32'hbcbb8cf5),
	.w3(32'hbc7fb31e),
	.w4(32'hbb5b738b),
	.w5(32'h3bf96d12),
	.w6(32'hbc7f9ad0),
	.w7(32'hbc374fd4),
	.w8(32'hbbc8d760),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb964be0),
	.w1(32'hbca5a363),
	.w2(32'hbb5d40a8),
	.w3(32'h39e4ec10),
	.w4(32'hbbda2eec),
	.w5(32'h3bd40de3),
	.w6(32'hbc2fc23e),
	.w7(32'h3bd6b3cb),
	.w8(32'h3c506d08),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b227b67),
	.w1(32'h3c4d7fed),
	.w2(32'hbcc84f98),
	.w3(32'hbbd97374),
	.w4(32'h3c83d117),
	.w5(32'h3ba95813),
	.w6(32'h3bb01e63),
	.w7(32'hbb9a44f1),
	.w8(32'h3c68bdad),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc40e31e),
	.w1(32'hbc91a6f3),
	.w2(32'hbc933615),
	.w3(32'hbcb66008),
	.w4(32'hbc95df8d),
	.w5(32'hbbcfb07a),
	.w6(32'h3c0684b1),
	.w7(32'hbc923363),
	.w8(32'h3caaa914),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca8604b),
	.w1(32'hbc0ef5fd),
	.w2(32'hbc056af4),
	.w3(32'h3cbf4322),
	.w4(32'hbb121c7a),
	.w5(32'hbc02ccd9),
	.w6(32'hbabdf9c1),
	.w7(32'hbc203de9),
	.w8(32'hb87489e1),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1e34d9),
	.w1(32'hbba7934f),
	.w2(32'hba5b8e85),
	.w3(32'h3af6c465),
	.w4(32'hbb2156bd),
	.w5(32'h3a102cb9),
	.w6(32'h3b6dd176),
	.w7(32'hb8a1d1c4),
	.w8(32'h3abf40fb),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba680ec),
	.w1(32'h3c616bbb),
	.w2(32'h3ab79d2c),
	.w3(32'h3b01b9cd),
	.w4(32'h3a02d347),
	.w5(32'hbc154d41),
	.w6(32'hbb459b36),
	.w7(32'hbbb5c153),
	.w8(32'h3a05559b),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae96830),
	.w1(32'hbb86d2a0),
	.w2(32'hbb984297),
	.w3(32'h3b44ab1e),
	.w4(32'hbb389588),
	.w5(32'hbbc99be1),
	.w6(32'hbb7ce73e),
	.w7(32'hbbfa7ee1),
	.w8(32'h3ccf82fa),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d20c001),
	.w1(32'hbc149794),
	.w2(32'hbc3063ff),
	.w3(32'h3d1164fb),
	.w4(32'hbb20ee38),
	.w5(32'hbb28c002),
	.w6(32'hbaad0ca0),
	.w7(32'hbbe62ca1),
	.w8(32'hbbae30b0),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbac5077),
	.w1(32'hbc238933),
	.w2(32'h3b824a94),
	.w3(32'hbb6e37cc),
	.w4(32'hbb9c5376),
	.w5(32'h3b6983f3),
	.w6(32'hbba65ed7),
	.w7(32'h3be74c70),
	.w8(32'hba0d4271),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7dd1a6),
	.w1(32'h3aaa7e3b),
	.w2(32'h3ba1e7a2),
	.w3(32'hbb535a2e),
	.w4(32'h3ab983c0),
	.w5(32'h3bbaefe3),
	.w6(32'h3b3a8793),
	.w7(32'h3c08d113),
	.w8(32'hbb49e8cc),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb58937f),
	.w1(32'hbb4eb173),
	.w2(32'hbb4c1ed6),
	.w3(32'hbb4fcbe5),
	.w4(32'hbb37aa0c),
	.w5(32'hbb51df18),
	.w6(32'hbb7b8698),
	.w7(32'hbb373b8e),
	.w8(32'h3b01da79),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb43720),
	.w1(32'hbbb83ca9),
	.w2(32'hbb99bbaf),
	.w3(32'h3ba213dd),
	.w4(32'hbbd0f869),
	.w5(32'hbbb57a68),
	.w6(32'hbb7f11b1),
	.w7(32'hbb7149fb),
	.w8(32'hbb2d2178),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb35a96a),
	.w1(32'hbb53726a),
	.w2(32'hbb252181),
	.w3(32'hbb48babc),
	.w4(32'hbb680434),
	.w5(32'hbb3eb591),
	.w6(32'hbb64ea25),
	.w7(32'hbb2f21d0),
	.w8(32'hbb621cc7),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb74f36f),
	.w1(32'hbb787c3e),
	.w2(32'hbb7691b5),
	.w3(32'hbb6bb79c),
	.w4(32'hbb7f939d),
	.w5(32'hbb8801bf),
	.w6(32'hbb70c9fa),
	.w7(32'hbb71606d),
	.w8(32'hbac62dae),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadc2691),
	.w1(32'hb9c4f957),
	.w2(32'hba0f8aba),
	.w3(32'hbb45e3d3),
	.w4(32'hbabe4c5a),
	.w5(32'hbaa547c7),
	.w6(32'hba0f6aec),
	.w7(32'hba2a1d0d),
	.w8(32'hbbafb3fe),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399b1513),
	.w1(32'hbb481805),
	.w2(32'hba0383b3),
	.w3(32'h3b1224b5),
	.w4(32'hba984780),
	.w5(32'hbadbf95a),
	.w6(32'hbb93bd39),
	.w7(32'h3a4849c3),
	.w8(32'hbb0ccc94),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4341ff),
	.w1(32'hba396967),
	.w2(32'hb9d09fa6),
	.w3(32'hbb3b0b18),
	.w4(32'hbac4e6f0),
	.w5(32'hba7f3421),
	.w6(32'hbabe0196),
	.w7(32'hbb13df71),
	.w8(32'h3bfe3e5a),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb8beb6),
	.w1(32'h3b912180),
	.w2(32'h3b835acd),
	.w3(32'h3c0678be),
	.w4(32'h3bf76689),
	.w5(32'h3bdd7ccd),
	.w6(32'h3bd49145),
	.w7(32'h3bc589b1),
	.w8(32'hbb61e047),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb572800),
	.w1(32'hbb4d5d87),
	.w2(32'hbb5c87e2),
	.w3(32'hbb5ef5c7),
	.w4(32'hbb4bcb16),
	.w5(32'hbb6f4b75),
	.w6(32'hbb5484de),
	.w7(32'hbb6a56c4),
	.w8(32'hbad9afec),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa68684),
	.w1(32'hba6d15d0),
	.w2(32'hba4f5f9d),
	.w3(32'hbaf152af),
	.w4(32'hbac7ed29),
	.w5(32'hbaaa6714),
	.w6(32'hbaaa1d4d),
	.w7(32'hba942661),
	.w8(32'hbb98e634),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb70d361),
	.w1(32'hbb3e06dd),
	.w2(32'hbb217495),
	.w3(32'hbb9855d4),
	.w4(32'hbb898379),
	.w5(32'hbb6560ba),
	.w6(32'hbb7ca608),
	.w7(32'hbb4a0359),
	.w8(32'hbb081957),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3ddfa8),
	.w1(32'h39d48c93),
	.w2(32'h3afff377),
	.w3(32'hbb2d35e5),
	.w4(32'hbb22ac7a),
	.w5(32'h3be4baa9),
	.w6(32'hbb77a2e4),
	.w7(32'h3b6c6319),
	.w8(32'h3b526c7c),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1a535e),
	.w1(32'hba18cd2b),
	.w2(32'hbacfb96b),
	.w3(32'h3b4617a7),
	.w4(32'h3b02f867),
	.w5(32'h3af7341f),
	.w6(32'hb991acac),
	.w7(32'hbadea1c4),
	.w8(32'hbbea7d8f),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb89e08),
	.w1(32'hbb29840b),
	.w2(32'hbb29e7b1),
	.w3(32'hbbc5c48c),
	.w4(32'hbb724a5f),
	.w5(32'hbb6be504),
	.w6(32'hbb70d1bb),
	.w7(32'hbba0de6e),
	.w8(32'h3ba68e5c),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb04b9f),
	.w1(32'hbb12ca89),
	.w2(32'hb9e946d8),
	.w3(32'hbb32bcc9),
	.w4(32'hbbd667ac),
	.w5(32'hb941efba),
	.w6(32'h3a5709ec),
	.w7(32'hbb300a7e),
	.w8(32'h3b0040b1),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b568d15),
	.w1(32'h3a7d6a57),
	.w2(32'h3a1e0130),
	.w3(32'h3b364904),
	.w4(32'hba31a479),
	.w5(32'hbb0f7d23),
	.w6(32'h3a865da1),
	.w7(32'h3975ee77),
	.w8(32'hbabb679b),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f7dff),
	.w1(32'hbb2c98c3),
	.w2(32'hbb618a12),
	.w3(32'hbba01fa7),
	.w4(32'hbb97ffc3),
	.w5(32'hbad1eafa),
	.w6(32'hbabfa0b6),
	.w7(32'hbba30737),
	.w8(32'h39f35960),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9c329d),
	.w1(32'hba6c8608),
	.w2(32'hbaba6768),
	.w3(32'h39f0594a),
	.w4(32'h3a9476f8),
	.w5(32'h39cddcbc),
	.w6(32'h3a41a50e),
	.w7(32'h3a5c713f),
	.w8(32'h3ab1f924),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a78e718),
	.w1(32'h392fc618),
	.w2(32'hbbc408d0),
	.w3(32'h3a7fa2e9),
	.w4(32'hbb769e22),
	.w5(32'hbba98a3a),
	.w6(32'hb9e089f0),
	.w7(32'hbbb0416d),
	.w8(32'hbb9013b4),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7e72f1),
	.w1(32'hba87bab6),
	.w2(32'hba0ad1cc),
	.w3(32'h3aa3dc67),
	.w4(32'hbba2ec39),
	.w5(32'hbb016e54),
	.w6(32'h37fecc8e),
	.w7(32'h3aaba411),
	.w8(32'hbac86cba),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba88f28c),
	.w1(32'hba3d3fe6),
	.w2(32'hbac606b1),
	.w3(32'hbb2bd5fa),
	.w4(32'hbb18ff9b),
	.w5(32'hbb0b9be3),
	.w6(32'hb97343bd),
	.w7(32'hba1d23be),
	.w8(32'hbba4569f),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba6f695),
	.w1(32'hbb662c09),
	.w2(32'hbb933b47),
	.w3(32'hbbba35f3),
	.w4(32'hbb86565d),
	.w5(32'hbba6893e),
	.w6(32'hbb8e422c),
	.w7(32'hbbb04f64),
	.w8(32'h39825377),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb95e06),
	.w1(32'hbb8e8d63),
	.w2(32'hbb858530),
	.w3(32'h3b38b56f),
	.w4(32'h3b42c526),
	.w5(32'h3adb0e46),
	.w6(32'hba8d5d51),
	.w7(32'hbb40d322),
	.w8(32'hbb00e01b),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule