module layer_10_featuremap_178(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3996c28b),
	.w1(32'h395e585b),
	.w2(32'hb7bb84aa),
	.w3(32'h39ba309e),
	.w4(32'h3a614cf1),
	.w5(32'h39aa35ee),
	.w6(32'hb9aa54ed),
	.w7(32'h38dafa1c),
	.w8(32'h3a20358b),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb35aa4f),
	.w1(32'hba1afc27),
	.w2(32'h3896790c),
	.w3(32'hbb4b90cc),
	.w4(32'h399cdb6b),
	.w5(32'h3aa58313),
	.w6(32'hbb46652f),
	.w7(32'hba93318d),
	.w8(32'h3a9dfe73),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38de1cfd),
	.w1(32'hb9b6cca5),
	.w2(32'hb9bcc658),
	.w3(32'hb84562a3),
	.w4(32'hb9b3a821),
	.w5(32'hb9a69c0c),
	.w6(32'hb81903c3),
	.w7(32'h378319b2),
	.w8(32'h389e976d),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3990e8a0),
	.w1(32'h3ac3533d),
	.w2(32'h3a67eed2),
	.w3(32'hb8c3b62a),
	.w4(32'h3aa9822d),
	.w5(32'h3a00fdc5),
	.w6(32'h3a0e989c),
	.w7(32'h39b1fb38),
	.w8(32'h3a8312f2),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95f0f90),
	.w1(32'h39a5c289),
	.w2(32'h39272bdf),
	.w3(32'hb977b045),
	.w4(32'h39dd45a6),
	.w5(32'h37ad31d0),
	.w6(32'h3915e07d),
	.w7(32'h388a279e),
	.w8(32'h38c0352b),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d8c82f),
	.w1(32'h3a127b0b),
	.w2(32'h3a2df688),
	.w3(32'h39b5e6f1),
	.w4(32'h39df3ede),
	.w5(32'h3a1bf075),
	.w6(32'h39e26c41),
	.w7(32'h39f3a732),
	.w8(32'h3a1bd297),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadb0b07),
	.w1(32'hbbfdfeaf),
	.w2(32'hbbae6206),
	.w3(32'h3b10399e),
	.w4(32'hbc1191b2),
	.w5(32'hbbbc9693),
	.w6(32'h3ad1db56),
	.w7(32'hbb6cb7ce),
	.w8(32'hbb200214),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb913c9b),
	.w1(32'hbb68494a),
	.w2(32'hbbabfb8c),
	.w3(32'hbb3fb79d),
	.w4(32'h3a966bb8),
	.w5(32'hbb822bde),
	.w6(32'h3b98c161),
	.w7(32'hbabb46b3),
	.w8(32'hbc5a1a0f),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2e03ac),
	.w1(32'hba328c3f),
	.w2(32'hba2e030a),
	.w3(32'hba4c31b3),
	.w4(32'hb8bdc4bc),
	.w5(32'hb9a4a81f),
	.w6(32'hba00965a),
	.w7(32'h3831e926),
	.w8(32'hba3cae34),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb101a33),
	.w1(32'hbac76d72),
	.w2(32'hbb4cae0f),
	.w3(32'h3a8e2b2f),
	.w4(32'h3abd5d01),
	.w5(32'h3a363d98),
	.w6(32'h3b6c43dc),
	.w7(32'h3ac1c9e8),
	.w8(32'h3aa96e5b),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b0921a),
	.w1(32'hb950c589),
	.w2(32'hb98ec8a3),
	.w3(32'hb9968705),
	.w4(32'hba557d7e),
	.w5(32'hba4cb46b),
	.w6(32'hb9ab004d),
	.w7(32'hb9e3c4f0),
	.w8(32'hba2158a3),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1149c9),
	.w1(32'hbb9f9f68),
	.w2(32'hbbad21bb),
	.w3(32'h3bab1ec4),
	.w4(32'hbb9a95c3),
	.w5(32'hbbfa694c),
	.w6(32'h3b9f8ef8),
	.w7(32'hbb318695),
	.w8(32'hbb04176e),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39823905),
	.w1(32'hbae93e71),
	.w2(32'hbb4daa51),
	.w3(32'h3b88596a),
	.w4(32'h3a6cfc0d),
	.w5(32'hb746bc82),
	.w6(32'h3bfa8bb6),
	.w7(32'h3b1d4eff),
	.w8(32'h389f0b08),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fef31a),
	.w1(32'hbb242bbc),
	.w2(32'hba6bc8f7),
	.w3(32'hb9adcf57),
	.w4(32'hbad89942),
	.w5(32'hba2d8fa6),
	.w6(32'hb92ab962),
	.w7(32'hbb0ebcc2),
	.w8(32'hba6862fc),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0cea12),
	.w1(32'h3a91ad51),
	.w2(32'h3b61cbaa),
	.w3(32'hbb485fd9),
	.w4(32'h3b1e3494),
	.w5(32'h3b632b2d),
	.w6(32'hbb260de6),
	.w7(32'h393994a0),
	.w8(32'h3b1a3a95),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a45b921),
	.w1(32'hb982bfbf),
	.w2(32'hbbce28ba),
	.w3(32'h3a6a2477),
	.w4(32'h3b8bb87d),
	.w5(32'h3a777dd5),
	.w6(32'hbac69de5),
	.w7(32'hbaecb28a),
	.w8(32'hbb8fa426),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8dd61ad),
	.w1(32'hb9b890e4),
	.w2(32'hb9dfbeec),
	.w3(32'hb8b9eed5),
	.w4(32'hba242639),
	.w5(32'hba4bfe1d),
	.w6(32'hba754fc2),
	.w7(32'hb9bf2d5d),
	.w8(32'hba1cebee),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab86cf5),
	.w1(32'hbbc70990),
	.w2(32'hbc2ddb2d),
	.w3(32'h3b7dc764),
	.w4(32'hbb926689),
	.w5(32'hbb9f4df1),
	.w6(32'h3bd60094),
	.w7(32'hb901000c),
	.w8(32'hbc351e98),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a151284),
	.w1(32'hbb3538b4),
	.w2(32'hbb8c3446),
	.w3(32'h3b7008c3),
	.w4(32'hba8b3a85),
	.w5(32'hbb1c7ef6),
	.w6(32'h3baf1921),
	.w7(32'h3ac457b9),
	.w8(32'hbb94c109),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb954c42d),
	.w1(32'h39948c20),
	.w2(32'h399dc163),
	.w3(32'hb9b2fe9f),
	.w4(32'h3a0a93d3),
	.w5(32'h39d335ef),
	.w6(32'hb954e97a),
	.w7(32'h3923b6f2),
	.w8(32'h38e4308d),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39416946),
	.w1(32'h39cabf86),
	.w2(32'h3979449c),
	.w3(32'h39df3506),
	.w4(32'h39f14841),
	.w5(32'h39acfaa3),
	.w6(32'h39eae5be),
	.w7(32'h39ae76bb),
	.w8(32'h38c2b03a),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1e8c28),
	.w1(32'h3a8b2c24),
	.w2(32'h3ad8bc1d),
	.w3(32'hb838f189),
	.w4(32'h3a963f91),
	.w5(32'h3ad5214e),
	.w6(32'hbb0e7ba4),
	.w7(32'hb7eea0ab),
	.w8(32'h3aaa7491),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc01b2cb),
	.w1(32'hbc176874),
	.w2(32'hbc8e76cd),
	.w3(32'h3a1552cc),
	.w4(32'hbba2d352),
	.w5(32'hbbcf5506),
	.w6(32'h3a6dde71),
	.w7(32'hbb7f5fd2),
	.w8(32'hba98c59c),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb63aa2b),
	.w1(32'hb9d43b87),
	.w2(32'h3a780ea2),
	.w3(32'hba8ed67d),
	.w4(32'h3b2d2670),
	.w5(32'h3b7e4c50),
	.w6(32'h3ac92553),
	.w7(32'h3b5a88ed),
	.w8(32'h3b9aeba0),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab4b4bd),
	.w1(32'h3b6d0a00),
	.w2(32'h3be3f07c),
	.w3(32'hbb10b9f7),
	.w4(32'h3bdd73de),
	.w5(32'h3c22e8a4),
	.w6(32'hbb971268),
	.w7(32'h3b8d3318),
	.w8(32'h3c125bbd),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c64cd2),
	.w1(32'hb9dbc359),
	.w2(32'hb9083d56),
	.w3(32'hb9d7799b),
	.w4(32'hb94cbd46),
	.w5(32'h36d2030f),
	.w6(32'hba16e408),
	.w7(32'hb986b7e7),
	.w8(32'h386b1349),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba72490b),
	.w1(32'h374fbc5d),
	.w2(32'h3933c85c),
	.w3(32'hba02a38e),
	.w4(32'h38f65d67),
	.w5(32'h395532f0),
	.w6(32'hb8ffdc20),
	.w7(32'hb8c12c22),
	.w8(32'hb956a3eb),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafd5349),
	.w1(32'hbade7d77),
	.w2(32'hbb6a0636),
	.w3(32'hba8d52ab),
	.w4(32'hbb7a5745),
	.w5(32'h3b4a20ad),
	.w6(32'hbb85b15a),
	.w7(32'hbba1a79a),
	.w8(32'h3a474695),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b75d01),
	.w1(32'hba7c8c5d),
	.w2(32'hb9ba0bbd),
	.w3(32'hb9d4edea),
	.w4(32'hba77ef0e),
	.w5(32'hb9a2bfba),
	.w6(32'h39080b69),
	.w7(32'hb805805c),
	.w8(32'h39b72b6b),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae96df9),
	.w1(32'h3b8e0dc0),
	.w2(32'h3c02f2f2),
	.w3(32'hbb213f5b),
	.w4(32'h3b3798be),
	.w5(32'h3c3d152d),
	.w6(32'hbba4a866),
	.w7(32'hbaf15c4b),
	.w8(32'h3c138d42),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39848503),
	.w1(32'h38a8819e),
	.w2(32'h382c68ca),
	.w3(32'hb8e75709),
	.w4(32'h3903628c),
	.w5(32'h390913b6),
	.w6(32'h38358683),
	.w7(32'h383b4b28),
	.w8(32'h366ed797),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb81ed04d),
	.w1(32'hb8bb1876),
	.w2(32'hb52adac2),
	.w3(32'h374f0fd2),
	.w4(32'hb6eb737b),
	.w5(32'h38f7c9f4),
	.w6(32'hb95507c9),
	.w7(32'hb90ba5de),
	.w8(32'hb9408e3f),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dd13e4),
	.w1(32'hb916fa80),
	.w2(32'hba1e8ab5),
	.w3(32'h3a9c8f39),
	.w4(32'h3a45eafb),
	.w5(32'h3a8dd525),
	.w6(32'h3accd02e),
	.w7(32'h3abe9fe0),
	.w8(32'h3a5f0631),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f88d5d),
	.w1(32'hba3c306e),
	.w2(32'h39eea9d2),
	.w3(32'hba8d3cde),
	.w4(32'h3a6198d3),
	.w5(32'h3a50d587),
	.w6(32'hbb336b35),
	.w7(32'hba2db8dc),
	.w8(32'hb90f5748),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a08042),
	.w1(32'hba248ad9),
	.w2(32'hba211b32),
	.w3(32'hb908a7d3),
	.w4(32'hb9941274),
	.w5(32'hba2e1919),
	.w6(32'hb951a329),
	.w7(32'hba2524f2),
	.w8(32'hba72d2b0),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb076abb),
	.w1(32'hbacecd0f),
	.w2(32'hbb3bca67),
	.w3(32'h3a62a297),
	.w4(32'hbad32562),
	.w5(32'hbb26f63b),
	.w6(32'h3b29538f),
	.w7(32'h39a47594),
	.w8(32'hb9c3c0b1),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc21ccd3),
	.w1(32'hbaa00b7f),
	.w2(32'hbc29cd70),
	.w3(32'hbc32752a),
	.w4(32'h3bbccb11),
	.w5(32'hbc407409),
	.w6(32'hbaa7c260),
	.w7(32'h3b23fef8),
	.w8(32'hb80e9546),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb70d6ac),
	.w1(32'h3c001ffa),
	.w2(32'h3c66e226),
	.w3(32'hbbde78bf),
	.w4(32'h3c06dea0),
	.w5(32'h3c8d71a0),
	.w6(32'hbbd0f950),
	.w7(32'h3be53bb7),
	.w8(32'h3c9e928d),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb54820),
	.w1(32'h3a32cab9),
	.w2(32'h3c43fa0b),
	.w3(32'hbbfdd2e1),
	.w4(32'hb732cd3b),
	.w5(32'h3c795e3d),
	.w6(32'hbbcad4c3),
	.w7(32'h3b81af35),
	.w8(32'h3c97249e),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399bac6e),
	.w1(32'h3adc4c97),
	.w2(32'h3b62b83f),
	.w3(32'h3a1ddacc),
	.w4(32'h3b2ca343),
	.w5(32'h3b499d40),
	.w6(32'hb91a4f0b),
	.w7(32'h3b0781e3),
	.w8(32'h3b3852bf),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e9cb23),
	.w1(32'hb980df85),
	.w2(32'hb9e3b4cd),
	.w3(32'hb9bb1c1c),
	.w4(32'hba0c1355),
	.w5(32'hba267d26),
	.w6(32'hb9c47bd2),
	.w7(32'hb9843ef5),
	.w8(32'hb9754cf7),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3999b8bc),
	.w1(32'h38e8b430),
	.w2(32'h39acf6c5),
	.w3(32'h3867d242),
	.w4(32'h38a69f13),
	.w5(32'h3946fa34),
	.w6(32'h396ea4b6),
	.w7(32'h39a500cc),
	.w8(32'h388c69a8),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cb00d7),
	.w1(32'hba651c25),
	.w2(32'hba09a1fd),
	.w3(32'hb982627f),
	.w4(32'hba45dedb),
	.w5(32'h37a0bdb4),
	.w6(32'hb9206918),
	.w7(32'hba357133),
	.w8(32'h39967c62),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad109a5),
	.w1(32'hbb341eb4),
	.w2(32'hbc2c0748),
	.w3(32'h3b32ae7d),
	.w4(32'h3a3e4d11),
	.w5(32'hbb6f9b19),
	.w6(32'h3bf970f7),
	.w7(32'h3ba5936a),
	.w8(32'hbb4e072a),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb161ebd),
	.w1(32'h3ab12246),
	.w2(32'h3b088365),
	.w3(32'hbafec9c9),
	.w4(32'h3b8b8d16),
	.w5(32'h3bc88c10),
	.w6(32'hbae508bb),
	.w7(32'h3b48f5a8),
	.w8(32'h3bc759e7),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb524c9a),
	.w1(32'hba3f5d35),
	.w2(32'h3afa0c9b),
	.w3(32'h383cfa65),
	.w4(32'h3b8db541),
	.w5(32'h3bbb2dab),
	.w6(32'h3adbfb8e),
	.w7(32'h3ba75456),
	.w8(32'h3bc22572),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9f14ed),
	.w1(32'hbaf294c9),
	.w2(32'hb9b49e9b),
	.w3(32'hbb661e10),
	.w4(32'h3acf8e98),
	.w5(32'h3a83454f),
	.w6(32'hb87aeb35),
	.w7(32'h3b0f013f),
	.w8(32'h3af1fc63),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb007e67),
	.w1(32'hbc237afb),
	.w2(32'hbc707f85),
	.w3(32'h3be26cd9),
	.w4(32'hbbb5a226),
	.w5(32'hbc093224),
	.w6(32'h3c37e25b),
	.w7(32'h3ad17de0),
	.w8(32'hbc13de7e),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cbf24b),
	.w1(32'hba1451da),
	.w2(32'hba43eb38),
	.w3(32'hba0be54b),
	.w4(32'hb8616aef),
	.w5(32'hb9f1724b),
	.w6(32'h37d3682f),
	.w7(32'h391575c0),
	.w8(32'hb93ab9c3),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ea279e),
	.w1(32'hb9cc267b),
	.w2(32'hb8a69667),
	.w3(32'h39b748c0),
	.w4(32'h3a499b26),
	.w5(32'h39809d3f),
	.w6(32'h39206d76),
	.w7(32'h3a25d907),
	.w8(32'hb8ae57d9),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3942e6a5),
	.w1(32'hb8a0696c),
	.w2(32'h35475a19),
	.w3(32'h39beaa1f),
	.w4(32'hb91afb2a),
	.w5(32'h3961a1b7),
	.w6(32'h3a77aaf4),
	.w7(32'h3a595ed4),
	.w8(32'h3a183f23),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb38d7d6),
	.w1(32'hba1e20eb),
	.w2(32'hbb033607),
	.w3(32'hba0063ce),
	.w4(32'h3a2e333c),
	.w5(32'h3abab6c5),
	.w6(32'hba2bfc7e),
	.w7(32'hb8917eda),
	.w8(32'h3b30bc61),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5ac91e),
	.w1(32'h38fe2292),
	.w2(32'hba03ce08),
	.w3(32'h3906b651),
	.w4(32'h39e6e901),
	.w5(32'h3831d995),
	.w6(32'h3ac6ab40),
	.w7(32'h3abf7d97),
	.w8(32'h39b8e33f),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a39e732),
	.w1(32'hbb8ce6eb),
	.w2(32'hbc0f5e8f),
	.w3(32'h3b9d9ea8),
	.w4(32'hbb0306dd),
	.w5(32'hbb942bdd),
	.w6(32'h3bf25616),
	.w7(32'hb91f7f14),
	.w8(32'hbc013ce2),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9aba431),
	.w1(32'hbb0ce87e),
	.w2(32'hbb3a8758),
	.w3(32'hba3e7ab9),
	.w4(32'hbb0d39e5),
	.w5(32'hbae6281a),
	.w6(32'hb9a24079),
	.w7(32'hb9a373c0),
	.w8(32'hbb0d6e72),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3917e4),
	.w1(32'h392ceb21),
	.w2(32'h39cef7dd),
	.w3(32'hba4e951f),
	.w4(32'h399f0d96),
	.w5(32'h39e0216f),
	.w6(32'h37d0c16c),
	.w7(32'h3994d98f),
	.w8(32'h3a1b0434),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e164a4),
	.w1(32'hb99621c0),
	.w2(32'hb9421dc7),
	.w3(32'h397e3aa0),
	.w4(32'hb98e4161),
	.w5(32'hb990378c),
	.w6(32'hb9a6c76b),
	.w7(32'h37fd2a93),
	.w8(32'h38a283c2),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90901b0),
	.w1(32'hb987bcb0),
	.w2(32'hb7090561),
	.w3(32'hb99b6d0a),
	.w4(32'hb9f73ffe),
	.w5(32'h3986d53f),
	.w6(32'hb9cc5d77),
	.w7(32'hb9e6b62f),
	.w8(32'h39882fca),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a00be45),
	.w1(32'h3a80d9d0),
	.w2(32'h3a8db896),
	.w3(32'hb930408a),
	.w4(32'h39f70408),
	.w5(32'h3a2bbeca),
	.w6(32'hb87217d8),
	.w7(32'h3a0217c5),
	.w8(32'h3a944fc8),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398bf4fa),
	.w1(32'hb8039307),
	.w2(32'h390a0cf0),
	.w3(32'hb8833623),
	.w4(32'hba061b2c),
	.w5(32'hb9bb3ac1),
	.w6(32'h390d26a7),
	.w7(32'hba1d1ed7),
	.w8(32'hba0bf6c2),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390caec0),
	.w1(32'hbb35f8b0),
	.w2(32'hbb981e7a),
	.w3(32'h3b0390c2),
	.w4(32'hbb04f8b3),
	.w5(32'hbb80aacb),
	.w6(32'h3b01163a),
	.w7(32'hb9bf0eb3),
	.w8(32'hbb9c4aa6),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f73cc9),
	.w1(32'hba6152f5),
	.w2(32'hbbeac012),
	.w3(32'hbb183268),
	.w4(32'hba741dab),
	.w5(32'hbb77890f),
	.w6(32'h3abbbeab),
	.w7(32'hba67b85e),
	.w8(32'hbbc8f5d5),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8959808),
	.w1(32'h3a2a59a5),
	.w2(32'h3945a5af),
	.w3(32'h39050c00),
	.w4(32'h3a94c6a4),
	.w5(32'h39ebbeea),
	.w6(32'h3689a0cc),
	.w7(32'h389b8190),
	.w8(32'h3916a17e),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8375471),
	.w1(32'h388eafd0),
	.w2(32'hb89380a3),
	.w3(32'hb91f11b8),
	.w4(32'hb941d415),
	.w5(32'hb985e0d7),
	.w6(32'h399b1352),
	.w7(32'h396cc7f9),
	.w8(32'h3a072ced),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39673ed5),
	.w1(32'hb9814aec),
	.w2(32'h38e606b0),
	.w3(32'hb861c953),
	.w4(32'hb9ea78e4),
	.w5(32'hb8ad8caf),
	.w6(32'hb8954cb2),
	.w7(32'hb7a27a48),
	.w8(32'h389a9008),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388426bc),
	.w1(32'hb9e26d7a),
	.w2(32'hba6c5053),
	.w3(32'h382ff769),
	.w4(32'hb9d709a7),
	.w5(32'hba27154a),
	.w6(32'hb9d48286),
	.w7(32'hba81db22),
	.w8(32'hba69218a),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395b7542),
	.w1(32'hbb9966c8),
	.w2(32'hbc101b6b),
	.w3(32'h3b02f522),
	.w4(32'hbaeb7b40),
	.w5(32'hbb80a9c3),
	.w6(32'h3bca211b),
	.w7(32'hbbd28e5c),
	.w8(32'hbc22d5f0),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa44751),
	.w1(32'hbb792c19),
	.w2(32'hbb3b9d6c),
	.w3(32'h3bc5d5d2),
	.w4(32'h3ad34a4a),
	.w5(32'hba1f3063),
	.w6(32'h3b04e15a),
	.w7(32'h3bbcf11d),
	.w8(32'hba201d4d),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcead4d),
	.w1(32'hbbbf2c8f),
	.w2(32'hbc1346b6),
	.w3(32'hbac422f8),
	.w4(32'hbb89c081),
	.w5(32'hbb97b761),
	.w6(32'h3aed692c),
	.w7(32'hba94326a),
	.w8(32'hbb8a8fad),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5f1e13),
	.w1(32'h3b9a4245),
	.w2(32'h3c137a20),
	.w3(32'hbbbc5346),
	.w4(32'h3bff97e8),
	.w5(32'h3c6afbb8),
	.w6(32'hbc0f531a),
	.w7(32'h3bd09b5e),
	.w8(32'h3c6b3d64),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb939baee),
	.w1(32'h394f4a8d),
	.w2(32'hb6e42974),
	.w3(32'hb9794dca),
	.w4(32'h3951efee),
	.w5(32'h382b2543),
	.w6(32'h393aee4c),
	.w7(32'h38ad7930),
	.w8(32'h39082edb),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3917d6eb),
	.w1(32'h390a1f5d),
	.w2(32'h37ffebd4),
	.w3(32'h37c68927),
	.w4(32'h388c3eb3),
	.w5(32'hb79ac985),
	.w6(32'h38137d71),
	.w7(32'h38a33005),
	.w8(32'hb8a63980),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394794b0),
	.w1(32'h39acf8db),
	.w2(32'h398e385a),
	.w3(32'h39652e01),
	.w4(32'h39b8c732),
	.w5(32'h3975f441),
	.w6(32'h395d0dcb),
	.w7(32'h39828f33),
	.w8(32'h39184905),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c35b80),
	.w1(32'hba93b8fa),
	.w2(32'hbb14b526),
	.w3(32'h3ab1b122),
	.w4(32'hb9fdd52a),
	.w5(32'hbae44dfe),
	.w6(32'h3b013733),
	.w7(32'h39ac1b6e),
	.w8(32'hbb377a9a),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392f534d),
	.w1(32'hb8d04ff6),
	.w2(32'hb8c4d150),
	.w3(32'h39ab53e6),
	.w4(32'hb7a39074),
	.w5(32'hb858c2b1),
	.w6(32'h397facd2),
	.w7(32'h39906eb9),
	.w8(32'h396fbdde),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad21d04),
	.w1(32'hbb68ed91),
	.w2(32'hbbd05917),
	.w3(32'h378c09ae),
	.w4(32'hbb1d2487),
	.w5(32'hbbb8b30c),
	.w6(32'h3b842b32),
	.w7(32'hbb06ce20),
	.w8(32'hbbad30ae),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1ecf20),
	.w1(32'hbaf9cd61),
	.w2(32'hbbadcc45),
	.w3(32'h3b703c7a),
	.w4(32'h38c742bc),
	.w5(32'hbbc99b32),
	.w6(32'h3bae951e),
	.w7(32'h3b15b497),
	.w8(32'hbbdebd17),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac978c2),
	.w1(32'h3a26573c),
	.w2(32'h3a888053),
	.w3(32'hbab64fd8),
	.w4(32'h3b84bfa1),
	.w5(32'h3b8033cf),
	.w6(32'hb93dcfe2),
	.w7(32'h3b22dab9),
	.w8(32'h3b68e2c1),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7311a8),
	.w1(32'hbb18af29),
	.w2(32'hbb8d4ed1),
	.w3(32'hba19e9bc),
	.w4(32'hbb295c58),
	.w5(32'hbb774272),
	.w6(32'h398a3c59),
	.w7(32'hbaf61084),
	.w8(32'hbbbd9a9a),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba37204a),
	.w1(32'hba07bd63),
	.w2(32'hba82d9b6),
	.w3(32'hba11c6db),
	.w4(32'h398c3d54),
	.w5(32'hba9f2a71),
	.w6(32'h3b067975),
	.w7(32'hbb0855bc),
	.w8(32'hbb73b066),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8c2dc0),
	.w1(32'hb963fa4c),
	.w2(32'hba90e3ea),
	.w3(32'hba94b3d7),
	.w4(32'h39b1a520),
	.w5(32'h3ab920ee),
	.w6(32'hba5857a7),
	.w7(32'h39bd48e3),
	.w8(32'h3a4b5b27),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba752b5f),
	.w1(32'hbb5eb33b),
	.w2(32'hbb976b90),
	.w3(32'h3ae0c0b7),
	.w4(32'hbb2ae4a1),
	.w5(32'hbb435cf0),
	.w6(32'h3b6d62bd),
	.w7(32'h39b1aa6e),
	.w8(32'hbb29e3f7),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39271a22),
	.w1(32'h39186398),
	.w2(32'h38324246),
	.w3(32'hb98c6752),
	.w4(32'h377d07ff),
	.w5(32'hb8445b3f),
	.w6(32'h39880bde),
	.w7(32'h39292a67),
	.w8(32'h39701ded),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3921c0df),
	.w1(32'hb981acb3),
	.w2(32'hb98aa46a),
	.w3(32'hb7d974d5),
	.w4(32'hb9c2ece6),
	.w5(32'hb9dc2536),
	.w6(32'hb93767d3),
	.w7(32'hb8074bf8),
	.w8(32'h38a9321b),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb69027ea),
	.w1(32'hba7897d5),
	.w2(32'hba33d925),
	.w3(32'hb92a511a),
	.w4(32'hba1d882b),
	.w5(32'hb9bc27bf),
	.w6(32'hba829c08),
	.w7(32'hba18ba13),
	.w8(32'hb9cabdf5),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa7071b),
	.w1(32'h39883b25),
	.w2(32'h3ae23d83),
	.w3(32'hbad73281),
	.w4(32'h38f446db),
	.w5(32'h3acd5231),
	.w6(32'hba3b0687),
	.w7(32'h39e77885),
	.w8(32'h3af8fd90),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaff84ad),
	.w1(32'hba016ba1),
	.w2(32'hba645ff9),
	.w3(32'hbb336883),
	.w4(32'h3b4c7b4d),
	.w5(32'h3a9a446a),
	.w6(32'hbb3d65f9),
	.w7(32'h3a9e2d37),
	.w8(32'h3b3972b9),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f391f6),
	.w1(32'h3a291777),
	.w2(32'h3a2c4b45),
	.w3(32'hba2224fd),
	.w4(32'h3a09e390),
	.w5(32'h3a439960),
	.w6(32'hb8b3d8ca),
	.w7(32'h395cbb58),
	.w8(32'h39d62f47),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3704d37b),
	.w1(32'hb96cd82f),
	.w2(32'h39e054f8),
	.w3(32'h3a219126),
	.w4(32'h3b355630),
	.w5(32'h3a35b403),
	.w6(32'hbaa670db),
	.w7(32'h3b04a09f),
	.w8(32'h39218cc4),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb045386),
	.w1(32'hbbc3a810),
	.w2(32'hbc0c1cd7),
	.w3(32'h3b12dea0),
	.w4(32'hbb7a773b),
	.w5(32'hbbc1e726),
	.w6(32'h3bb58db6),
	.w7(32'h3881d52d),
	.w8(32'hbc0a7ad2),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5e4a7c),
	.w1(32'hba05617e),
	.w2(32'h3b5d7541),
	.w3(32'hbb802447),
	.w4(32'h3931b63b),
	.w5(32'h3bc01541),
	.w6(32'hbb311ca6),
	.w7(32'h3b2fbb36),
	.w8(32'h3c14e07d),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0c01bb),
	.w1(32'hbb00d735),
	.w2(32'hbc1609d2),
	.w3(32'h3b88d73c),
	.w4(32'h3aa7bb64),
	.w5(32'hbb9e5830),
	.w6(32'h3aa4ad79),
	.w7(32'hbaacd7ff),
	.w8(32'h3a46b74b),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90004c1),
	.w1(32'h3b0dbd2a),
	.w2(32'h3b9311d1),
	.w3(32'hbaee2dd4),
	.w4(32'h3b5dedf6),
	.w5(32'h3bbb6891),
	.w6(32'h3a01768d),
	.w7(32'h3bb71be6),
	.w8(32'h3c021f91),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac6f154),
	.w1(32'hbaef3df4),
	.w2(32'hbb8efb8f),
	.w3(32'h3a92c53d),
	.w4(32'h3996b8e2),
	.w5(32'hbaa12f0a),
	.w6(32'h3a35cebf),
	.w7(32'hba5fa82c),
	.w8(32'hbbe7c7e8),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba89bf2f),
	.w1(32'hbaeb0bc9),
	.w2(32'hbb076f43),
	.w3(32'hbae3ea2e),
	.w4(32'hba3a3ccb),
	.w5(32'hba44ae87),
	.w6(32'hbb02c806),
	.w7(32'hbb323da0),
	.w8(32'hbb0eb81a),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafd591d),
	.w1(32'h3b86eff6),
	.w2(32'h3bf66d31),
	.w3(32'hbb59c243),
	.w4(32'h3b997954),
	.w5(32'h3c10af39),
	.w6(32'hbb701515),
	.w7(32'h3b2586b1),
	.w8(32'h3c0f53dc),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa162aa),
	.w1(32'hba661a92),
	.w2(32'hbaa39226),
	.w3(32'h3a2a1471),
	.w4(32'hba779c30),
	.w5(32'hba0d38b2),
	.w6(32'hba3a0e71),
	.w7(32'hba6cff9d),
	.w8(32'hba19b7d9),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac90514),
	.w1(32'hbac84ba5),
	.w2(32'hbb6000fa),
	.w3(32'h3b0c12a5),
	.w4(32'h3a9e58fc),
	.w5(32'h3a4bfab1),
	.w6(32'h3ba59104),
	.w7(32'h3b524375),
	.w8(32'hba944a7d),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9601c87),
	.w1(32'hbbbe7ae1),
	.w2(32'hbbd84851),
	.w3(32'h3a36c8a1),
	.w4(32'hbb0879c0),
	.w5(32'hbb28440f),
	.w6(32'h3bc217eb),
	.w7(32'h3956e303),
	.w8(32'h3b0084aa),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc65d2aa),
	.w1(32'hba20057f),
	.w2(32'hbc333821),
	.w3(32'h3b830370),
	.w4(32'h3c009bd6),
	.w5(32'hbc1f7d36),
	.w6(32'h3b2b5aea),
	.w7(32'h3b83cdb5),
	.w8(32'h3abe8d9a),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb28c919),
	.w1(32'h3b5c96e7),
	.w2(32'h3c19180c),
	.w3(32'hbba86e2e),
	.w4(32'h3c061739),
	.w5(32'h3c63e9be),
	.w6(32'hbbc7efeb),
	.w7(32'h3c1a4c48),
	.w8(32'h3cacac11),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f10d12),
	.w1(32'h3b4af7ba),
	.w2(32'h3bb0fceb),
	.w3(32'hb9dd67c8),
	.w4(32'h3bd6fbdb),
	.w5(32'h3c0e6873),
	.w6(32'hba10c1a1),
	.w7(32'h3bb74b92),
	.w8(32'h3bf11e37),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeb9522),
	.w1(32'hbb9bf8ab),
	.w2(32'hbc294e4d),
	.w3(32'h3a5394b4),
	.w4(32'h38b9ac17),
	.w5(32'hbc0e2aff),
	.w6(32'h3ae6f13b),
	.w7(32'hbb279ced),
	.w8(32'hba75952d),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac071d3),
	.w1(32'hba392f60),
	.w2(32'hbae42e57),
	.w3(32'h3ab3e40b),
	.w4(32'hb8759889),
	.w5(32'hb9ed750d),
	.w6(32'h3a5c763c),
	.w7(32'h38b75ff2),
	.w8(32'h3806786f),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3e685d),
	.w1(32'hbbcc95c0),
	.w2(32'hbc3e7083),
	.w3(32'hbbf2ab1d),
	.w4(32'h3b6641ba),
	.w5(32'hbc4958bc),
	.w6(32'hbc06884a),
	.w7(32'hbb79ded0),
	.w8(32'hbb807af8),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb59ef87),
	.w1(32'hbab319c1),
	.w2(32'hbb77bdd4),
	.w3(32'hb8be39f0),
	.w4(32'h3b0b5608),
	.w5(32'hbb846dce),
	.w6(32'h3bc0ed9c),
	.w7(32'h3abbe083),
	.w8(32'h3a884ef1),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89fee89),
	.w1(32'hba0ba8b8),
	.w2(32'hb9e1d329),
	.w3(32'hb804095f),
	.w4(32'hba27ec2b),
	.w5(32'hb9db2a56),
	.w6(32'hba2252ff),
	.w7(32'hb9bf6a51),
	.w8(32'h38d44780),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabba0b6),
	.w1(32'hbaa7f028),
	.w2(32'hbb1447ef),
	.w3(32'h398ab844),
	.w4(32'h3a816ba3),
	.w5(32'h3963f379),
	.w6(32'hbaaeffe7),
	.w7(32'hba058819),
	.w8(32'h3990a6c2),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3591269c),
	.w1(32'hba796c3f),
	.w2(32'hbb3d34c8),
	.w3(32'h3b5487d1),
	.w4(32'h3afe84cd),
	.w5(32'h3abf8da2),
	.w6(32'h3bc1255a),
	.w7(32'h3b7026e9),
	.w8(32'h3a9e0f03),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacb384b),
	.w1(32'h3b078671),
	.w2(32'h3b8ff700),
	.w3(32'hba5620fb),
	.w4(32'h3b9c8a92),
	.w5(32'h3be772c0),
	.w6(32'hba3be810),
	.w7(32'h3b81e9e8),
	.w8(32'h3bda70a1),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9fffb8),
	.w1(32'hba77bccf),
	.w2(32'h3b07234b),
	.w3(32'hbb8439cc),
	.w4(32'h3a6fb0b7),
	.w5(32'h3bc4e502),
	.w6(32'hbade4928),
	.w7(32'h3afff8eb),
	.w8(32'h3c02e0f2),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1b056f),
	.w1(32'hb91cba6f),
	.w2(32'h39c3426c),
	.w3(32'hbb3e81f8),
	.w4(32'h3b5947d7),
	.w5(32'h3b46513c),
	.w6(32'hbb200734),
	.w7(32'h3a096cfb),
	.w8(32'h3b2c09de),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8513f2),
	.w1(32'h3b4d6d6f),
	.w2(32'h3ae94ad0),
	.w3(32'h3b51fc83),
	.w4(32'h3b62e078),
	.w5(32'h3a4cd36b),
	.w6(32'h3ac8dfe6),
	.w7(32'h3b3fb9bf),
	.w8(32'hb98ab5b2),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a93cae),
	.w1(32'hbb4bc012),
	.w2(32'hbbd38fc7),
	.w3(32'hb951e0e7),
	.w4(32'hba8a17c8),
	.w5(32'hbb6855ec),
	.w6(32'hbb05720c),
	.w7(32'hbb8a5cbd),
	.w8(32'hbb9838bd),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba951bdc),
	.w1(32'hb978007c),
	.w2(32'h3a1493bc),
	.w3(32'hba7cd4bb),
	.w4(32'h3ab8781c),
	.w5(32'h3b1e5fc5),
	.w6(32'hb9d822cb),
	.w7(32'h3a916ecc),
	.w8(32'h3b1e46af),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6b9ad9),
	.w1(32'hb90c88f4),
	.w2(32'hb99c25c3),
	.w3(32'hba6275f6),
	.w4(32'hb8ab8bfb),
	.w5(32'hb9714f47),
	.w6(32'hb9a83e6a),
	.w7(32'hb95cba84),
	.w8(32'h3840bc13),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb81cf329),
	.w1(32'hb8a9f12b),
	.w2(32'hba6b0e48),
	.w3(32'hb92687d4),
	.w4(32'h390a768e),
	.w5(32'hba32e7d1),
	.w6(32'hb973ca4c),
	.w7(32'hba75c626),
	.w8(32'hbaadbedf),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399718f5),
	.w1(32'h3992dbb7),
	.w2(32'h395e0d21),
	.w3(32'h398fb9eb),
	.w4(32'h398f2ad8),
	.w5(32'h3982c41d),
	.w6(32'h3928ca62),
	.w7(32'h393a5c38),
	.w8(32'h3977fe82),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c31289),
	.w1(32'h38eaf655),
	.w2(32'hb9de6a22),
	.w3(32'h39a1ed8f),
	.w4(32'h39e98ca1),
	.w5(32'h38cfd2d2),
	.w6(32'hba2db3b7),
	.w7(32'hb94b3a3c),
	.w8(32'hb98615d1),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba929470),
	.w1(32'h3a989d86),
	.w2(32'h3b1c13d6),
	.w3(32'hba1b8933),
	.w4(32'h3b51d996),
	.w5(32'h3b942196),
	.w6(32'h39a8d2a6),
	.w7(32'h3b45fbea),
	.w8(32'h3b78a071),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39721841),
	.w1(32'hb8b83c68),
	.w2(32'hba5ee78d),
	.w3(32'h39898eff),
	.w4(32'hb85c9a70),
	.w5(32'hb9fcd033),
	.w6(32'hb9264b11),
	.w7(32'h3930d93c),
	.w8(32'hb9a4a841),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb926bd31),
	.w1(32'hb983a56c),
	.w2(32'hbb33b4ad),
	.w3(32'h3b01badc),
	.w4(32'hb982012e),
	.w5(32'hbafe0ee1),
	.w6(32'h3b561229),
	.w7(32'h3a7152e8),
	.w8(32'hbab4a854),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4422d7),
	.w1(32'h3af46edb),
	.w2(32'h3bab7886),
	.w3(32'hbb584e35),
	.w4(32'h3b6c812e),
	.w5(32'h3c074266),
	.w6(32'hbb940b78),
	.w7(32'h3aa317a1),
	.w8(32'h3bfeea04),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39249b06),
	.w1(32'hb9cbeb3a),
	.w2(32'hba24c632),
	.w3(32'h3932cf9c),
	.w4(32'hb9303105),
	.w5(32'hb976d704),
	.w6(32'hba663749),
	.w7(32'hb85291ee),
	.w8(32'hb7966c5d),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dba760),
	.w1(32'h3a123b28),
	.w2(32'h3a097e38),
	.w3(32'hba0a50f6),
	.w4(32'h3a0af9b4),
	.w5(32'h39dc009d),
	.w6(32'h3a499872),
	.w7(32'h3a4c2da1),
	.w8(32'h3a2d2fa9),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8b4bbe),
	.w1(32'h39454c44),
	.w2(32'h394af798),
	.w3(32'h3a7b4a04),
	.w4(32'h3965f1ec),
	.w5(32'h396096c9),
	.w6(32'h3975302f),
	.w7(32'h39196286),
	.w8(32'h38a9fa4d),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb84914d0),
	.w1(32'hb8b987d0),
	.w2(32'hbb001406),
	.w3(32'h39ee7474),
	.w4(32'h3a802239),
	.w5(32'hba9110ba),
	.w6(32'h3aad86ef),
	.w7(32'hbaafb352),
	.w8(32'h39f5850b),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad2b728),
	.w1(32'hbb690b1a),
	.w2(32'hbb8a76a4),
	.w3(32'h3b934288),
	.w4(32'hbb851a2f),
	.w5(32'hbb5d7aa3),
	.w6(32'h3b65c4d4),
	.w7(32'h3b38acb3),
	.w8(32'hbb1fbec2),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb996adfa),
	.w1(32'hb8252d4d),
	.w2(32'hbbc95a26),
	.w3(32'h3b5f9301),
	.w4(32'h3b17ff63),
	.w5(32'hbadd4c11),
	.w6(32'h3ba9f366),
	.w7(32'hba2aef1e),
	.w8(32'hbb9ef1b6),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a30cdbb),
	.w1(32'hbb01d520),
	.w2(32'hbb4dbc4b),
	.w3(32'h39ec165a),
	.w4(32'hba89a8b6),
	.w5(32'hbafda459),
	.w6(32'hbab45bff),
	.w7(32'hbb1b9345),
	.w8(32'hbb031151),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbace92ab),
	.w1(32'hbb3c77be),
	.w2(32'hbb191938),
	.w3(32'hb9a8de65),
	.w4(32'hbab974c0),
	.w5(32'hbb1fb826),
	.w6(32'hbb025c61),
	.w7(32'hbad3fffc),
	.w8(32'hbb93f210),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1169f2),
	.w1(32'hbab0a76f),
	.w2(32'hb9c44a6b),
	.w3(32'hbab0ab2f),
	.w4(32'h3ade7cd9),
	.w5(32'h3af93dc2),
	.w6(32'h3a94b125),
	.w7(32'h3a56df5b),
	.w8(32'h3b0cbfd5),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadd66e4),
	.w1(32'h392b0b2d),
	.w2(32'hbad97f0d),
	.w3(32'h398be056),
	.w4(32'hba174c59),
	.w5(32'h3ac00a1d),
	.w6(32'h3a48baac),
	.w7(32'h3aa3add1),
	.w8(32'hbaa0b695),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa8c1f4),
	.w1(32'hbb95fb17),
	.w2(32'hbba93a8f),
	.w3(32'hbaa30c53),
	.w4(32'hbb2a0d0c),
	.w5(32'hbae65469),
	.w6(32'hbb3ef712),
	.w7(32'hbb822242),
	.w8(32'hbb955421),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad44e43),
	.w1(32'hbbf47e61),
	.w2(32'hbc37d9ac),
	.w3(32'h3b55faac),
	.w4(32'hbbe549ba),
	.w5(32'hbbd3b9dd),
	.w6(32'h3af1b78c),
	.w7(32'hbb971ab8),
	.w8(32'hbbf900b8),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafe7db9),
	.w1(32'h3b0e2235),
	.w2(32'h3ace5da2),
	.w3(32'hbb246311),
	.w4(32'h3b6f9904),
	.w5(32'h3b59b2fd),
	.w6(32'hbb624009),
	.w7(32'h3ad384c9),
	.w8(32'h3b55605f),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafedf38),
	.w1(32'hbac916e7),
	.w2(32'hbb28bd01),
	.w3(32'h3ad886b1),
	.w4(32'h3a5def93),
	.w5(32'h39ad7e5d),
	.w6(32'h3ac09e91),
	.w7(32'h3b23679f),
	.w8(32'h3a9ebfa0),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9abc12),
	.w1(32'hbb93bf92),
	.w2(32'hbbc56161),
	.w3(32'h3b680570),
	.w4(32'hbb2534c7),
	.w5(32'hbab5a439),
	.w6(32'h3b7037d2),
	.w7(32'hba1d0ae2),
	.w8(32'hba4668ae),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abf5375),
	.w1(32'hb9edf485),
	.w2(32'hba3b3c95),
	.w3(32'h3b981ed4),
	.w4(32'h3b7bb91f),
	.w5(32'h3a7b7164),
	.w6(32'hba367e9a),
	.w7(32'h3b80928f),
	.w8(32'h3aeeb691),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9b1226),
	.w1(32'h3a53a004),
	.w2(32'hba2fca99),
	.w3(32'h3a790c08),
	.w4(32'hba1df01c),
	.w5(32'hbb017c93),
	.w6(32'h3b03b828),
	.w7(32'hb93b906e),
	.w8(32'hb909e4ae),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb940a312),
	.w1(32'h398cd6ae),
	.w2(32'hba1b70f7),
	.w3(32'hba68f0c2),
	.w4(32'h3acf429f),
	.w5(32'h3a382362),
	.w6(32'h3a575b29),
	.w7(32'h38825aa8),
	.w8(32'h39f872b0),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a042e46),
	.w1(32'h3bc1cf96),
	.w2(32'h3c2f6fa7),
	.w3(32'hbb164281),
	.w4(32'h3bac352b),
	.w5(32'h3c5432c7),
	.w6(32'hbc0e5194),
	.w7(32'h39fe8471),
	.w8(32'h3c33788b),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8db101),
	.w1(32'h3afdcecd),
	.w2(32'h3ab76b03),
	.w3(32'hbb4abcbd),
	.w4(32'hba10e37e),
	.w5(32'h3a0284d0),
	.w6(32'h3acc6bf9),
	.w7(32'h3b5fa69a),
	.w8(32'h3b1a37a4),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b36a45e),
	.w1(32'h39e1a3da),
	.w2(32'h37c081cb),
	.w3(32'h3b1f5d8a),
	.w4(32'h39146e1c),
	.w5(32'h38fe2f4f),
	.w6(32'hb8a69612),
	.w7(32'h375eba2d),
	.w8(32'hba2280c1),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38acc1bb),
	.w1(32'h38fac9ee),
	.w2(32'h3a20de73),
	.w3(32'hb9d95c45),
	.w4(32'hba3c2e56),
	.w5(32'hb7317968),
	.w6(32'h3a82b567),
	.w7(32'h3b3e7dbd),
	.w8(32'hba1a22ee),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb196b8b),
	.w1(32'hb9fc4279),
	.w2(32'hba5cacfe),
	.w3(32'h382e3555),
	.w4(32'h39b954ff),
	.w5(32'h388adfb4),
	.w6(32'hbae38050),
	.w7(32'hba14d9d3),
	.w8(32'h3aa9d794),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5ad326),
	.w1(32'h38069916),
	.w2(32'h38493f91),
	.w3(32'hbb0add3f),
	.w4(32'h3b56f34a),
	.w5(32'h3b2d77ac),
	.w6(32'hbb4da10f),
	.w7(32'h3a28f845),
	.w8(32'h3b171473),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaad17b5),
	.w1(32'hbab670ec),
	.w2(32'hba8d1f44),
	.w3(32'h3b67d6f0),
	.w4(32'h3ae636aa),
	.w5(32'h3ad3e9da),
	.w6(32'h3bb84608),
	.w7(32'h3b83b1d4),
	.w8(32'h399cf1e2),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399b07fa),
	.w1(32'h3a5a754e),
	.w2(32'hb9de2d9d),
	.w3(32'h380eb79d),
	.w4(32'h3aa2c825),
	.w5(32'hba2b2c5a),
	.w6(32'h3aead9c3),
	.w7(32'hb96d38c0),
	.w8(32'hb9e1acbe),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb05b8dc),
	.w1(32'hba584609),
	.w2(32'hbb07465d),
	.w3(32'hba504dd0),
	.w4(32'h3a7c6b03),
	.w5(32'hb8a699cf),
	.w6(32'h3b768563),
	.w7(32'h39a18c37),
	.w8(32'hbb72c927),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb20c1da),
	.w1(32'h3b55727b),
	.w2(32'h39c87561),
	.w3(32'hbaa8f55a),
	.w4(32'h3bd263ce),
	.w5(32'h3b37c0d4),
	.w6(32'h3be7eeab),
	.w7(32'h3b4d0576),
	.w8(32'h3b495ef4),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0e4e29),
	.w1(32'hbb9102b9),
	.w2(32'hbc0c0aa8),
	.w3(32'h3b25f215),
	.w4(32'hbaceb274),
	.w5(32'hbb91c32b),
	.w6(32'h3b016283),
	.w7(32'hbae28f85),
	.w8(32'hbb58f9ec),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbc0a71),
	.w1(32'h3ac663e9),
	.w2(32'h389244fb),
	.w3(32'hbb91a43c),
	.w4(32'h3a1eb8dd),
	.w5(32'h3be1b348),
	.w6(32'hbb1373cd),
	.w7(32'hba47378a),
	.w8(32'h3bc25fa1),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7af404),
	.w1(32'hbb158dfe),
	.w2(32'hb8c8ee38),
	.w3(32'hba293647),
	.w4(32'hbafb68eb),
	.w5(32'hba85dfdb),
	.w6(32'hbad13478),
	.w7(32'hbac1914b),
	.w8(32'h3a012b09),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5973f6),
	.w1(32'h3ad8d690),
	.w2(32'h3a1cc7ac),
	.w3(32'h3b142b66),
	.w4(32'h3b1ed17b),
	.w5(32'h3aafb2a6),
	.w6(32'h3ae15bad),
	.w7(32'h3ab9f867),
	.w8(32'h3acafc73),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba10a47a),
	.w1(32'h3b06c0f9),
	.w2(32'h3a28323a),
	.w3(32'hbab99c0f),
	.w4(32'h3b7711f7),
	.w5(32'h3ba92a0d),
	.w6(32'hbab8f537),
	.w7(32'h3af89297),
	.w8(32'h3b9ac3ae),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1c9f6a),
	.w1(32'hbad3d9ca),
	.w2(32'h3b241c8f),
	.w3(32'hbadbc285),
	.w4(32'h3a626e7a),
	.w5(32'h3bc14ddf),
	.w6(32'hba9ed2f3),
	.w7(32'h3bdbbb88),
	.w8(32'h3ae2c31c),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb615f3f),
	.w1(32'h3b10499a),
	.w2(32'h3acef48a),
	.w3(32'hbb3478e0),
	.w4(32'h3a2e7b77),
	.w5(32'h3b080451),
	.w6(32'h39e25a64),
	.w7(32'h3a503557),
	.w8(32'h3a4733c9),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1b6f5d),
	.w1(32'hb96c2bf9),
	.w2(32'hbb1f7bea),
	.w3(32'hbae6e19f),
	.w4(32'h392a58d8),
	.w5(32'hbaea9711),
	.w6(32'h3adc590f),
	.w7(32'hba7f41f9),
	.w8(32'hba97aac0),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c1ab8b),
	.w1(32'hb994aa16),
	.w2(32'hba802a85),
	.w3(32'hb78ff159),
	.w4(32'h3a526dd7),
	.w5(32'hba1cf68c),
	.w6(32'h39a45c65),
	.w7(32'hbaa8566c),
	.w8(32'hb9bde7ab),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97fef26),
	.w1(32'hb99599f3),
	.w2(32'hbb32ea6e),
	.w3(32'h3b1b6dd1),
	.w4(32'h399e5390),
	.w5(32'h3a79e529),
	.w6(32'h3b60cbfd),
	.w7(32'h3b0fc014),
	.w8(32'hba1b09c0),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a29f789),
	.w1(32'h3bcaaf0c),
	.w2(32'hbbf18f0e),
	.w3(32'h3a950b39),
	.w4(32'h3c469579),
	.w5(32'hbbb9b757),
	.w6(32'h3c30eebd),
	.w7(32'hbba6d834),
	.w8(32'h3b44bed0),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b270ffa),
	.w1(32'h3a3a1ca1),
	.w2(32'hb98dc9fe),
	.w3(32'h3947a372),
	.w4(32'h3abf47e4),
	.w5(32'h3b707e35),
	.w6(32'hbb9b2cea),
	.w7(32'hbac721a4),
	.w8(32'h3afc67cf),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba12546e),
	.w1(32'h3a88f6a4),
	.w2(32'h39cadc42),
	.w3(32'h3a4217cc),
	.w4(32'h3a581845),
	.w5(32'h39ae58a0),
	.w6(32'h3a793f40),
	.w7(32'hb8ab9a2e),
	.w8(32'h396f7d0e),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb955a6f3),
	.w1(32'hbb132f33),
	.w2(32'hb7c35e27),
	.w3(32'h3a9d58d3),
	.w4(32'hbb5d08dc),
	.w5(32'hb9eef22d),
	.w6(32'hbae15a51),
	.w7(32'hbab0e4a2),
	.w8(32'hbaf7f931),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb963cff5),
	.w1(32'hba816c18),
	.w2(32'hbb061798),
	.w3(32'h3a9939fb),
	.w4(32'hba6c4889),
	.w5(32'hbabc163d),
	.w6(32'hbabdd3ab),
	.w7(32'hbaf844d8),
	.w8(32'hba584a31),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f5925b),
	.w1(32'hba6a2c43),
	.w2(32'hbac7b0d6),
	.w3(32'h392db353),
	.w4(32'hba34cfd5),
	.w5(32'hbaa1c5a9),
	.w6(32'hba8af6bd),
	.w7(32'hba86c44f),
	.w8(32'hba695155),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb67234a),
	.w1(32'hba6261a6),
	.w2(32'hbab7514f),
	.w3(32'hbb94be1e),
	.w4(32'hb97a3a18),
	.w5(32'h3a984a31),
	.w6(32'hbba6e528),
	.w7(32'hbaeda795),
	.w8(32'h3a53d9cf),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb993128),
	.w1(32'h3ae61365),
	.w2(32'hbbe19bec),
	.w3(32'h3b1fc018),
	.w4(32'h3bb29698),
	.w5(32'hbb2f5f95),
	.w6(32'h3c464504),
	.w7(32'h3b85bb60),
	.w8(32'hbaddd5cd),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb255fa8),
	.w1(32'hb8108227),
	.w2(32'hb96757b6),
	.w3(32'hbb4675c1),
	.w4(32'hba52a7c9),
	.w5(32'hb9e49a9d),
	.w6(32'hba748026),
	.w7(32'hba20f1fd),
	.w8(32'hb97d3c59),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0d6cbc),
	.w1(32'h3b148541),
	.w2(32'h3b7d29ac),
	.w3(32'hbb17cba3),
	.w4(32'h3bb45ec2),
	.w5(32'h3bc6bb64),
	.w6(32'h39468a52),
	.w7(32'h3b036efd),
	.w8(32'h3b977817),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a92f2ad),
	.w1(32'hbb22ddfe),
	.w2(32'hbb0aa461),
	.w3(32'h3ac44997),
	.w4(32'hba9532dd),
	.w5(32'h3b0bd709),
	.w6(32'hba002b2a),
	.w7(32'h3a3235c7),
	.w8(32'h3af2f6c2),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b08958c),
	.w1(32'hbba7b653),
	.w2(32'hbc1ec27b),
	.w3(32'h3b9b94b0),
	.w4(32'hbb37e150),
	.w5(32'hbba42579),
	.w6(32'h399d0660),
	.w7(32'hb9d40079),
	.w8(32'hbbe63cf5),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb52362b),
	.w1(32'hbb9580e5),
	.w2(32'hbbb7dce3),
	.w3(32'hba8bed2e),
	.w4(32'hbaba6ab4),
	.w5(32'hbaae4fa4),
	.w6(32'hb81b5f0a),
	.w7(32'hbaf49d8a),
	.w8(32'hbaba0b5a),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb189950),
	.w1(32'hb90e727e),
	.w2(32'hbb5ebed1),
	.w3(32'hba41eaf1),
	.w4(32'hbae12b43),
	.w5(32'hbb3297e5),
	.w6(32'h3ba06cdf),
	.w7(32'h3b43a74c),
	.w8(32'hbabacb28),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acecfdf),
	.w1(32'h3ad44ef7),
	.w2(32'h3ad434e3),
	.w3(32'h3a63e2d4),
	.w4(32'h3b72403a),
	.w5(32'h3b81d3c4),
	.w6(32'h3bc4a3b8),
	.w7(32'h3bf161da),
	.w8(32'h3a2fcd9a),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb532e39),
	.w1(32'hb9b08262),
	.w2(32'hbaf4fa16),
	.w3(32'hbb1c0dc8),
	.w4(32'h3aa3e7ac),
	.w5(32'hba7950bb),
	.w6(32'h38821c5f),
	.w7(32'hbae4d2fa),
	.w8(32'hbb35549a),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a21d791),
	.w1(32'hba408224),
	.w2(32'hba98cc02),
	.w3(32'h3a402a0d),
	.w4(32'hba67e3e9),
	.w5(32'hba394b43),
	.w6(32'hba844138),
	.w7(32'hba35cba1),
	.w8(32'hba56b18d),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac69fee),
	.w1(32'hbb0467a6),
	.w2(32'hbb41e1a5),
	.w3(32'hba8e7d88),
	.w4(32'hbb2b4087),
	.w5(32'hbb1e7c05),
	.w6(32'hbb0e16a3),
	.w7(32'hbabd67be),
	.w8(32'hb9000c6d),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac1750b),
	.w1(32'h3ba37c8d),
	.w2(32'hbbc4aae2),
	.w3(32'hbb0c7c10),
	.w4(32'h3b1e3768),
	.w5(32'h390f4a38),
	.w6(32'h3b23f239),
	.w7(32'hbaee534f),
	.w8(32'h3847c06e),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabdb55a),
	.w1(32'h3a2999ba),
	.w2(32'hbb059531),
	.w3(32'hb9a0b6f2),
	.w4(32'h3b3b45c1),
	.w5(32'h3a327066),
	.w6(32'h3a21d2b7),
	.w7(32'h383b22d8),
	.w8(32'hbaf8c618),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7aa84c),
	.w1(32'hba858705),
	.w2(32'h3af4eca4),
	.w3(32'h398f5b2e),
	.w4(32'hbaac05bf),
	.w5(32'h3ad1d09c),
	.w6(32'hb8b9276d),
	.w7(32'h3add23f2),
	.w8(32'h398bc5c3),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c5f202),
	.w1(32'hbad24534),
	.w2(32'hbaaa7f70),
	.w3(32'h3a34f54c),
	.w4(32'hba393ccd),
	.w5(32'hb9dac800),
	.w6(32'hba067f62),
	.w7(32'hb9f13991),
	.w8(32'hb92030a4),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9b8173),
	.w1(32'hba686865),
	.w2(32'h39dfa49e),
	.w3(32'hb9fa860e),
	.w4(32'hbac26e9c),
	.w5(32'h3add8670),
	.w6(32'hbb427de0),
	.w7(32'hba73a9f6),
	.w8(32'hba9607b6),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc05ee8b),
	.w1(32'hbba6fae5),
	.w2(32'hbbfff572),
	.w3(32'hbba7d2a5),
	.w4(32'hbaceedd1),
	.w5(32'hbbbe3511),
	.w6(32'hbb00b29f),
	.w7(32'hbba11abb),
	.w8(32'hbb65eb4c),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc10fdd0),
	.w1(32'h3b45be6f),
	.w2(32'hbc31ebc9),
	.w3(32'hbbe9520e),
	.w4(32'h3b8c7c9a),
	.w5(32'hbbc66adb),
	.w6(32'h3a8435c7),
	.w7(32'hbacc43a2),
	.w8(32'hbb06aa17),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba99c1e5),
	.w1(32'hbb09f386),
	.w2(32'hbb94fbdb),
	.w3(32'hba5aa751),
	.w4(32'hbabd7276),
	.w5(32'hbb3a1ae5),
	.w6(32'hbb36ec07),
	.w7(32'hbb74ce14),
	.w8(32'hbb48d543),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a84960f),
	.w1(32'hbb07c987),
	.w2(32'hbbd0a8fb),
	.w3(32'h3bf1e5bd),
	.w4(32'h39ae322b),
	.w5(32'hbb9dc5ca),
	.w6(32'h3c248fa0),
	.w7(32'h3b0a5edd),
	.w8(32'hbbdf1a78),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf1abb8),
	.w1(32'hb96c7367),
	.w2(32'hbbf4a248),
	.w3(32'hbbfd19f3),
	.w4(32'h3a87090b),
	.w5(32'h3aafca7e),
	.w6(32'hbb825374),
	.w7(32'hbb5cfdab),
	.w8(32'h3a17f476),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba179d94),
	.w1(32'hbab6e3a2),
	.w2(32'hbaf70556),
	.w3(32'hb9c896bb),
	.w4(32'hba391048),
	.w5(32'hbad7a42f),
	.w6(32'h3a0770ff),
	.w7(32'h384f1a29),
	.w8(32'hbb58cf0d),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba901122),
	.w1(32'h3a1563d0),
	.w2(32'hbb0b5cf7),
	.w3(32'hb9575ed2),
	.w4(32'hb97c863b),
	.w5(32'hb917373c),
	.w6(32'hba299481),
	.w7(32'hbb3c3163),
	.w8(32'hbb1be56d),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafab490),
	.w1(32'hbad71282),
	.w2(32'h39df2031),
	.w3(32'hbae13672),
	.w4(32'hb9914878),
	.w5(32'h3b04898c),
	.w6(32'hbaad5ddd),
	.w7(32'h3a664831),
	.w8(32'h3b0ec702),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ada7a93),
	.w1(32'hba838f27),
	.w2(32'hba2b4886),
	.w3(32'h3b328502),
	.w4(32'hba830037),
	.w5(32'h39927f6e),
	.w6(32'hba526ff5),
	.w7(32'hb8f0292b),
	.w8(32'hba440d2f),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac01d5a),
	.w1(32'hbabb616c),
	.w2(32'hbc064484),
	.w3(32'h3abc4b07),
	.w4(32'hbb0fb4c8),
	.w5(32'hbb85f333),
	.w6(32'h3a3b4ce1),
	.w7(32'hbb40778f),
	.w8(32'hb87cccec),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadb7c85),
	.w1(32'h3b2d5f96),
	.w2(32'hbab1e858),
	.w3(32'h3a49f0f6),
	.w4(32'h3ab557f3),
	.w5(32'hbb1214af),
	.w6(32'h3bd72c47),
	.w7(32'h39c364a0),
	.w8(32'hb9f376cd),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa091eb),
	.w1(32'h3bbfc43c),
	.w2(32'hbb38e2ca),
	.w3(32'hbb142d92),
	.w4(32'h3c3ca513),
	.w5(32'hb9db4c76),
	.w6(32'h3c30cc41),
	.w7(32'hb93f4d2b),
	.w8(32'h3a46bdae),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb71d87d),
	.w1(32'h3a50d12c),
	.w2(32'h3a816504),
	.w3(32'hbb14d3ae),
	.w4(32'h3a3aa632),
	.w5(32'h3a27415e),
	.w6(32'hba0dd337),
	.w7(32'h3a366663),
	.w8(32'h3a79d723),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadf85c0),
	.w1(32'hbb996287),
	.w2(32'hbc18dbbe),
	.w3(32'h3aa74990),
	.w4(32'hbb3fbdd5),
	.w5(32'hbb73d8b5),
	.w6(32'h3a9363dc),
	.w7(32'hbacab759),
	.w8(32'hba3a373f),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb90266b),
	.w1(32'hbb0f3482),
	.w2(32'hbb7357fa),
	.w3(32'hbb0dd45c),
	.w4(32'h394cb4b1),
	.w5(32'hbb4e5308),
	.w6(32'hbadca109),
	.w7(32'hbad20c97),
	.w8(32'hbaaab567),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb906992d),
	.w1(32'h3826adce),
	.w2(32'hbaa52baa),
	.w3(32'h39b8bee6),
	.w4(32'hb9100c2d),
	.w5(32'hba8fd1a3),
	.w6(32'hba054667),
	.w7(32'hba839725),
	.w8(32'hba95e7f9),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0f40dc),
	.w1(32'hba2d3e5b),
	.w2(32'hbb79c9fb),
	.w3(32'hbaa67774),
	.w4(32'h3a2f5342),
	.w5(32'hbb06b629),
	.w6(32'hbae04d52),
	.w7(32'hbabd9f25),
	.w8(32'hbb1ec31b),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8200b9),
	.w1(32'h3a30d213),
	.w2(32'hb9fe6fb2),
	.w3(32'hba3096cb),
	.w4(32'h3aa4f60c),
	.w5(32'hb9bce45f),
	.w6(32'h3a99eb83),
	.w7(32'hba42b4bf),
	.w8(32'hb8dd6e42),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb49835e),
	.w1(32'hbb8b0ab2),
	.w2(32'hbbc0de7e),
	.w3(32'h39bd87ab),
	.w4(32'hbb231ef2),
	.w5(32'hbaaace0a),
	.w6(32'hba4b0da3),
	.w7(32'hbaf0f69e),
	.w8(32'hbb036e9e),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb88b2a1),
	.w1(32'h3aa8495b),
	.w2(32'h3b616976),
	.w3(32'hbb89a8bb),
	.w4(32'h3ab94574),
	.w5(32'h3ac98434),
	.w6(32'hbb4de449),
	.w7(32'h3a50a5e9),
	.w8(32'h3baa5bd1),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba116d54),
	.w1(32'hba8b4699),
	.w2(32'h3a58bab6),
	.w3(32'hba962ee9),
	.w4(32'h3acb5797),
	.w5(32'h3b7056f9),
	.w6(32'hbac9e633),
	.w7(32'h3b06d7f7),
	.w8(32'h3b84a3d0),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a4cffe),
	.w1(32'hba3e2f15),
	.w2(32'hbb08875a),
	.w3(32'h3a4a8d4a),
	.w4(32'hbac28e85),
	.w5(32'hba889a4f),
	.w6(32'hbaf8d189),
	.w7(32'hbb062219),
	.w8(32'hbae25a70),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9269d1),
	.w1(32'hba49a5f2),
	.w2(32'h3a81d24c),
	.w3(32'hbb96d044),
	.w4(32'h3b1c4ceb),
	.w5(32'h3bb4d930),
	.w6(32'hbb76c623),
	.w7(32'h3ab64084),
	.w8(32'h3b835fda),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2e1ba4),
	.w1(32'h3ac3c8df),
	.w2(32'hbaf5f1dc),
	.w3(32'h3b787433),
	.w4(32'h3b488b53),
	.w5(32'h3a200a7b),
	.w6(32'h3b3c2065),
	.w7(32'h39dff512),
	.w8(32'hb9ffc213),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba18dd3a),
	.w1(32'h3c0228b5),
	.w2(32'hbb7db0ce),
	.w3(32'h3b6d74c4),
	.w4(32'h3c43ff4b),
	.w5(32'hbb4eeb3d),
	.w6(32'h3c997fa5),
	.w7(32'h3a2a54bd),
	.w8(32'hba57ce43),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1f399b),
	.w1(32'hb9dec141),
	.w2(32'hba849dd9),
	.w3(32'hbb1324cd),
	.w4(32'hba9a4a5e),
	.w5(32'hbae1c8ff),
	.w6(32'hba6e8775),
	.w7(32'hbaa5ba5e),
	.w8(32'hbaf2ce27),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae58c71),
	.w1(32'h3a3f77d6),
	.w2(32'h3a10a664),
	.w3(32'hbb0d0aec),
	.w4(32'hb815ba62),
	.w5(32'h39773072),
	.w6(32'h3a4f0f7e),
	.w7(32'h3a79c3e3),
	.w8(32'hb9aee4bc),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb95f2fe),
	.w1(32'hbb7c60c1),
	.w2(32'hbbdaee4d),
	.w3(32'h3a747e60),
	.w4(32'hb63abb48),
	.w5(32'hbb8fb916),
	.w6(32'h3a92825e),
	.w7(32'h3a7f1845),
	.w8(32'hbb31a691),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba75933),
	.w1(32'h3b13644a),
	.w2(32'hbc156757),
	.w3(32'h39ae63e7),
	.w4(32'h3c226ef6),
	.w5(32'hbbbd7815),
	.w6(32'h3c536b28),
	.w7(32'h39b0ccbe),
	.w8(32'h3b019952),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb92e959),
	.w1(32'h3afe277b),
	.w2(32'h3b3a5cd5),
	.w3(32'hbac7ce48),
	.w4(32'h3b7e21c3),
	.w5(32'h3b9a52ed),
	.w6(32'h3aae4a52),
	.w7(32'h3b62f8dc),
	.w8(32'h3b38669d),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5c3f08),
	.w1(32'hbba33e73),
	.w2(32'hbb90b910),
	.w3(32'hbaeb87d1),
	.w4(32'hbbae38cc),
	.w5(32'hbb684612),
	.w6(32'h39b031e1),
	.w7(32'hbbb7f22a),
	.w8(32'hbb9cbc22),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf781bd),
	.w1(32'h3aa9065c),
	.w2(32'h3a29b0e1),
	.w3(32'hbaf5c5bb),
	.w4(32'h3aa9115b),
	.w5(32'h3a28eb03),
	.w6(32'h3a88b9e4),
	.w7(32'h39f653ea),
	.w8(32'h397e0f74),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88b3140),
	.w1(32'hba51e2b1),
	.w2(32'hbb067a7f),
	.w3(32'h3a194cbe),
	.w4(32'hb9b37c1e),
	.w5(32'hbaa9d83a),
	.w6(32'h39a09dd3),
	.w7(32'hba83bfa8),
	.w8(32'hbac96b43),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ed944),
	.w1(32'hb9270288),
	.w2(32'hbc0f1232),
	.w3(32'h3b92b6d0),
	.w4(32'h3b132f9c),
	.w5(32'hbbd6db89),
	.w6(32'h3bed616c),
	.w7(32'h3b80d80d),
	.w8(32'h3bc7115d),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaf6438),
	.w1(32'hbb3ac8b5),
	.w2(32'hbbb7d8cb),
	.w3(32'h3bdc6240),
	.w4(32'hba32a9f8),
	.w5(32'hbb9976db),
	.w6(32'h3c09e5f2),
	.w7(32'h3a8354eb),
	.w8(32'hbbba820a),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba2a09b),
	.w1(32'hbb12f4dc),
	.w2(32'hbc037eb6),
	.w3(32'h3b565269),
	.w4(32'h3a3fea09),
	.w5(32'hbbcf548a),
	.w6(32'h3b3a6640),
	.w7(32'h3b1c1f64),
	.w8(32'h391c60c7),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e7373e),
	.w1(32'h3b0a09f1),
	.w2(32'h3b77bb24),
	.w3(32'hba46f311),
	.w4(32'h3b3ef5d9),
	.w5(32'h3bb0d354),
	.w6(32'hbaeea155),
	.w7(32'h3b101e8d),
	.w8(32'h3bab3145),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb897ff3),
	.w1(32'h3ba1646b),
	.w2(32'h3aa30089),
	.w3(32'hbb9cd4fb),
	.w4(32'h3bfb4fb2),
	.w5(32'h3b9e8f3f),
	.w6(32'h3ad209be),
	.w7(32'hba4d3bd1),
	.w8(32'h3b47e694),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb332257),
	.w1(32'hba9e5b98),
	.w2(32'hbace2c25),
	.w3(32'hbb28b7f6),
	.w4(32'hba2586f5),
	.w5(32'hba17612b),
	.w6(32'hbac583d1),
	.w7(32'hbaad134a),
	.w8(32'hba97a9f8),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8da78a),
	.w1(32'hb963eac8),
	.w2(32'h3aed230b),
	.w3(32'hba10fba3),
	.w4(32'h39e046d4),
	.w5(32'h39ee9449),
	.w6(32'h39e0269c),
	.w7(32'h3afb0c35),
	.w8(32'h3a58dc3b),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9233448),
	.w1(32'h3bfcd2cc),
	.w2(32'hbb4601a1),
	.w3(32'hba3c576b),
	.w4(32'h3bfe0582),
	.w5(32'hbb37ffa1),
	.w6(32'h3c32b361),
	.w7(32'hbafee2e6),
	.w8(32'hbad58437),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba80727b),
	.w1(32'h3aaefeac),
	.w2(32'hbb2825e9),
	.w3(32'hb99c8e81),
	.w4(32'h3b07afbd),
	.w5(32'h3b0bc0e1),
	.w6(32'h3ab6958f),
	.w7(32'hb8c08fc3),
	.w8(32'hb973c676),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba017da6),
	.w1(32'hbb7e3a60),
	.w2(32'hbb84d065),
	.w3(32'hb94d41ff),
	.w4(32'hbb855315),
	.w5(32'hbb6711c7),
	.w6(32'hba5f0db3),
	.w7(32'hbba006ef),
	.w8(32'hbb3bac4d),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab3f21d),
	.w1(32'h3ab824ad),
	.w2(32'h398d06a9),
	.w3(32'h3b19b04e),
	.w4(32'h3b2cdb70),
	.w5(32'h3af334df),
	.w6(32'h3ac93afb),
	.w7(32'h3b4560ed),
	.w8(32'h3a7048d2),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac4889b),
	.w1(32'hbac06333),
	.w2(32'hbbbc630d),
	.w3(32'h37ecea31),
	.w4(32'h391dab68),
	.w5(32'hba05754d),
	.w6(32'hba822ad8),
	.w7(32'hba9744d3),
	.w8(32'h3b294eda),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d6e122),
	.w1(32'h3b158331),
	.w2(32'hbac62df6),
	.w3(32'hbacfb96a),
	.w4(32'h3b4135f1),
	.w5(32'h39fd6b92),
	.w6(32'h3aecb948),
	.w7(32'hb8a7d62e),
	.w8(32'h3a4b910a),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb96b078),
	.w1(32'hbb7f0f8c),
	.w2(32'hbc29e62e),
	.w3(32'h3b60e5fc),
	.w4(32'hb9d97baa),
	.w5(32'hbba437d7),
	.w6(32'h3b4565a8),
	.w7(32'h3ba9d007),
	.w8(32'hba6f13cb),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fd67e1),
	.w1(32'hbaad16b6),
	.w2(32'hbb742daa),
	.w3(32'h3b6dc7db),
	.w4(32'hba85fde2),
	.w5(32'hbb45fc6d),
	.w6(32'h3a735560),
	.w7(32'hbaad283f),
	.w8(32'hbb654a09),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba989cbd),
	.w1(32'hba83fb28),
	.w2(32'hb9892236),
	.w3(32'hbabca376),
	.w4(32'hb9aa873f),
	.w5(32'h3a399eb3),
	.w6(32'hba5e9b19),
	.w7(32'h39c31185),
	.w8(32'h3a214585),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8a8ce7),
	.w1(32'hb94f9461),
	.w2(32'hbad3f74b),
	.w3(32'h3b9b698e),
	.w4(32'h3a9cf472),
	.w5(32'h399d894b),
	.w6(32'h3b964aa0),
	.w7(32'h3b340335),
	.w8(32'hb8b01bff),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9b78a3),
	.w1(32'hbaf9f70d),
	.w2(32'hbad01ed1),
	.w3(32'h3a9327d0),
	.w4(32'hba91a5ce),
	.w5(32'hba4174d1),
	.w6(32'hbb24d9f0),
	.w7(32'hbb13bcaf),
	.w8(32'hbb15a7ff),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadab185),
	.w1(32'h3a9fdca5),
	.w2(32'hb8af0269),
	.w3(32'hb9f13be6),
	.w4(32'h3acc8717),
	.w5(32'hb9dd1901),
	.w6(32'h3b164827),
	.w7(32'h39a16611),
	.w8(32'hb8f076c9),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8f290b),
	.w1(32'hba554f9b),
	.w2(32'hb9c2eb60),
	.w3(32'hba7ef732),
	.w4(32'hb89d42e9),
	.w5(32'h3a0a82ed),
	.w6(32'hba2adeb1),
	.w7(32'h39ef7ea5),
	.w8(32'h39ffc8bf),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8dedf29),
	.w1(32'hbb88a19d),
	.w2(32'hbb8669ab),
	.w3(32'h3a433ffc),
	.w4(32'hbb8af7dc),
	.w5(32'hbb6de623),
	.w6(32'hbb901843),
	.w7(32'hbb946b4f),
	.w8(32'hbb83620b),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5f6fb0),
	.w1(32'h3a85866f),
	.w2(32'hba039078),
	.w3(32'hbb710c7e),
	.w4(32'h39e360fd),
	.w5(32'h375598ba),
	.w6(32'hba9f37d9),
	.w7(32'hba539198),
	.w8(32'h3a9f8960),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb37bc82),
	.w1(32'hbba58af9),
	.w2(32'hbbdd1349),
	.w3(32'hba7a3abe),
	.w4(32'hba72bfdc),
	.w5(32'h3b13e120),
	.w6(32'h3aac795c),
	.w7(32'hbb569a05),
	.w8(32'hbb94f5a4),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39807517),
	.w1(32'hba807815),
	.w2(32'hbb76ac14),
	.w3(32'h3b2cff52),
	.w4(32'hb963c514),
	.w5(32'hbab136b1),
	.w6(32'h3af69bb7),
	.w7(32'h3a6f8fc4),
	.w8(32'hbac5a8eb),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab1fa20),
	.w1(32'hbba7b4fd),
	.w2(32'hbc16d079),
	.w3(32'h3a74cdba),
	.w4(32'hbb95a8ad),
	.w5(32'hbbb78a1a),
	.w6(32'h3a51ba8d),
	.w7(32'hbb80b6cc),
	.w8(32'hbbdacf57),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2cab27),
	.w1(32'hba643735),
	.w2(32'h3a8b96f0),
	.w3(32'hbb03848a),
	.w4(32'h39e2d064),
	.w5(32'h3a8d79a0),
	.w6(32'hb98ffe2f),
	.w7(32'hba5587cf),
	.w8(32'hba2c7180),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a46f7ee),
	.w1(32'hbaac2617),
	.w2(32'hb9bce740),
	.w3(32'h3a3ba1ba),
	.w4(32'hb9885f4b),
	.w5(32'h3a456e66),
	.w6(32'hba2a5e3a),
	.w7(32'h3a1c994f),
	.w8(32'h3980a150),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88c3875),
	.w1(32'hba151a54),
	.w2(32'hba516575),
	.w3(32'h3aa6a675),
	.w4(32'hb946815c),
	.w5(32'hb9725fe4),
	.w6(32'hba172e8f),
	.w7(32'hb8fd0a3a),
	.w8(32'hb9c18211),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba56eef3),
	.w1(32'hba43573a),
	.w2(32'hb96bcb4e),
	.w3(32'hb851ae69),
	.w4(32'hb97180ec),
	.w5(32'h3a2bfad1),
	.w6(32'hba61e3ae),
	.w7(32'h3a23bdd4),
	.w8(32'h38be7bf2),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8557f5),
	.w1(32'hbb451830),
	.w2(32'hbb9468d1),
	.w3(32'h3a0abbca),
	.w4(32'hba84ec28),
	.w5(32'hbb6f249a),
	.w6(32'h38ceefa1),
	.w7(32'h3a4fbe88),
	.w8(32'hbbfc7fb2),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae63696),
	.w1(32'hbaa0c0be),
	.w2(32'hbabcfbcd),
	.w3(32'hba886791),
	.w4(32'hbac4b5f8),
	.w5(32'h3aa7afb7),
	.w6(32'hba9c4da4),
	.w7(32'h3ab4e8a9),
	.w8(32'hba0ec798),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fbf64c),
	.w1(32'h3aa91203),
	.w2(32'h3a6d8349),
	.w3(32'h37a2c9ed),
	.w4(32'h3ae1a26e),
	.w5(32'h3a42785c),
	.w6(32'h3aa1a6d6),
	.w7(32'h38d334e1),
	.w8(32'h39d5f4a3),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9f972f),
	.w1(32'h3b06a14a),
	.w2(32'h39d5322f),
	.w3(32'h39371158),
	.w4(32'h3b35be0b),
	.w5(32'h3aab75c0),
	.w6(32'h3a5480a7),
	.w7(32'h3add1273),
	.w8(32'hb999fb3d),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397c6d70),
	.w1(32'hbab0326f),
	.w2(32'hbaf86e1e),
	.w3(32'h3a094524),
	.w4(32'hba6e0281),
	.w5(32'hbab584e9),
	.w6(32'hbaaa8e80),
	.w7(32'hba9cd1a7),
	.w8(32'hbab5f33c),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb22e373),
	.w1(32'hb95bb36b),
	.w2(32'h3a641419),
	.w3(32'hb99fceec),
	.w4(32'h3b080064),
	.w5(32'hba2a1b44),
	.w6(32'h3b79eda0),
	.w7(32'h3b3868d7),
	.w8(32'hb96adf32),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99c58f9),
	.w1(32'h3a2f5310),
	.w2(32'h3b2ae952),
	.w3(32'h39c00ff3),
	.w4(32'h3aa992e0),
	.w5(32'h3ad41b72),
	.w6(32'h39959bbc),
	.w7(32'h3ab8f219),
	.w8(32'h3a066d7a),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a995404),
	.w1(32'hbb436a8c),
	.w2(32'hbc52b6a7),
	.w3(32'h3b1288a4),
	.w4(32'h3adca078),
	.w5(32'hbb9b405b),
	.w6(32'h3b1a47d2),
	.w7(32'hbab8769f),
	.w8(32'hbc140d35),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3765fcf8),
	.w1(32'h3c032a25),
	.w2(32'hbad85a9c),
	.w3(32'hb85cb194),
	.w4(32'hbc057029),
	.w5(32'h3c0cbe20),
	.w6(32'hbc00ca33),
	.w7(32'h3a90b313),
	.w8(32'h3bf545e6),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ec1ade),
	.w1(32'h3d197488),
	.w2(32'h3b53a2d9),
	.w3(32'h3c4ba5ec),
	.w4(32'h3c314dd5),
	.w5(32'h3beeba0c),
	.w6(32'h3bc6571a),
	.w7(32'h3b7b8cb6),
	.w8(32'hbbc74445),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule