module layer_8_featuremap_28(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9be4816),
	.w1(32'hba2e21ed),
	.w2(32'h38e58f55),
	.w3(32'hba4ea133),
	.w4(32'hba773d47),
	.w5(32'hb98b92a7),
	.w6(32'h39df897c),
	.w7(32'h39cc1c2f),
	.w8(32'h3a1939e0),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2cb441),
	.w1(32'h39a4bdef),
	.w2(32'h3a504396),
	.w3(32'h3b2fdb1a),
	.w4(32'h3a1ba9c3),
	.w5(32'h3a5d629b),
	.w6(32'h3b4d92ab),
	.w7(32'h3adb545e),
	.w8(32'h3b2a50ee),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9dfd05),
	.w1(32'h3aa04245),
	.w2(32'h3b3acb2c),
	.w3(32'h3baab188),
	.w4(32'h3afed35f),
	.w5(32'h3b1d12de),
	.w6(32'h3bc1d632),
	.w7(32'h3b194f18),
	.w8(32'h3b3fb75f),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba51b313),
	.w1(32'hb895233d),
	.w2(32'h3ae451d1),
	.w3(32'hba508a2a),
	.w4(32'hbab94271),
	.w5(32'hb9d88e5d),
	.w6(32'h39b80c2c),
	.w7(32'hb9847bfb),
	.w8(32'h39e9d952),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b871c65),
	.w1(32'h3b533f45),
	.w2(32'h3ba8f3bb),
	.w3(32'h3b7d4def),
	.w4(32'h3b3533a9),
	.w5(32'h3ba43e8d),
	.w6(32'h3ba8285c),
	.w7(32'h3b8b8fa7),
	.w8(32'h3c06e4ca),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2ad070),
	.w1(32'hbb43293f),
	.w2(32'h3b2b0c38),
	.w3(32'h3b9371c7),
	.w4(32'hbb0426e9),
	.w5(32'h3b097e43),
	.w6(32'h3b16208c),
	.w7(32'h3b158689),
	.w8(32'h3a1dd977),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9792055),
	.w1(32'hba1a48af),
	.w2(32'hba0f3849),
	.w3(32'hb969be66),
	.w4(32'hb9e3aa19),
	.w5(32'hba55226f),
	.w6(32'hba2b2e35),
	.w7(32'hba38eaf4),
	.w8(32'h39e91f47),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2b29b9),
	.w1(32'h3a58e119),
	.w2(32'h3abf3d53),
	.w3(32'h3aff2389),
	.w4(32'hba10636a),
	.w5(32'h3ae20cd5),
	.w6(32'h3b69e859),
	.w7(32'h3b1faaa3),
	.w8(32'h3b3e2239),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4c7f7d),
	.w1(32'h3a8f86a4),
	.w2(32'h3b3c26cf),
	.w3(32'h3b51bd20),
	.w4(32'h3ae02b0a),
	.w5(32'h3aeb81d8),
	.w6(32'h3ba5999f),
	.w7(32'h3b0bb931),
	.w8(32'h3b934e2a),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b434497),
	.w1(32'h3b31535e),
	.w2(32'h3b961ca5),
	.w3(32'hb9d2ed5e),
	.w4(32'hbb66c3e7),
	.w5(32'hba01de9b),
	.w6(32'h3baa6710),
	.w7(32'h3b199ae8),
	.w8(32'h3b26097d),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf41dcc),
	.w1(32'h392ab996),
	.w2(32'h3b00d751),
	.w3(32'hbb3cd0db),
	.w4(32'hba676e49),
	.w5(32'h3a935ab8),
	.w6(32'hbb3824dd),
	.w7(32'hba8d6823),
	.w8(32'hba95faaa),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8cdc13d),
	.w1(32'hba554bbd),
	.w2(32'h37fcb86e),
	.w3(32'hb9daeb28),
	.w4(32'hba51a066),
	.w5(32'hba5cfdb9),
	.w6(32'hb7859fd5),
	.w7(32'hb9c0bcc7),
	.w8(32'h3a84f96d),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0ac7a4),
	.w1(32'hba363809),
	.w2(32'h3a886d80),
	.w3(32'h3b311021),
	.w4(32'hb8a6bd82),
	.w5(32'h39d703c7),
	.w6(32'h3b6968b5),
	.w7(32'h3a40722b),
	.w8(32'h3bee313d),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b277efc),
	.w1(32'hbb39e9f4),
	.w2(32'h3a5c120e),
	.w3(32'h3bb1eb78),
	.w4(32'hba039122),
	.w5(32'h3afc3393),
	.w6(32'h3ab0d80b),
	.w7(32'h3b6bca50),
	.w8(32'h398e2f65),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a784f9f),
	.w1(32'hb9d04ee0),
	.w2(32'h3a87de79),
	.w3(32'h3b00bac2),
	.w4(32'h389abb27),
	.w5(32'h39f0a63c),
	.w6(32'h3a85b3a2),
	.w7(32'h3abcc91d),
	.w8(32'h399e8ed4),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4002d7),
	.w1(32'h3a2017b1),
	.w2(32'h3a053e0a),
	.w3(32'h390fd992),
	.w4(32'h392abe61),
	.w5(32'h38818ca4),
	.w6(32'h3987a9df),
	.w7(32'h39203816),
	.w8(32'h3ab0fe17),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3ad120),
	.w1(32'hbb0704a9),
	.w2(32'h3a7785cd),
	.w3(32'h3af604bb),
	.w4(32'h3b647baa),
	.w5(32'h3bdb5bdb),
	.w6(32'h3a26b064),
	.w7(32'h3a5dc186),
	.w8(32'h3ae1675b),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b69f2fd),
	.w1(32'h3a3fb9ae),
	.w2(32'h3b021c38),
	.w3(32'h3b6cb0a4),
	.w4(32'h3a554abe),
	.w5(32'h3ab3ae21),
	.w6(32'h3b8f44b8),
	.w7(32'h3b26abb0),
	.w8(32'h3b430ac2),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2022eb),
	.w1(32'hbab19fd3),
	.w2(32'h3bbf34b9),
	.w3(32'hbb876619),
	.w4(32'hbb90dbfb),
	.w5(32'h3b399c9a),
	.w6(32'hbaf55df5),
	.w7(32'hbb7b07b0),
	.w8(32'h3b54ea4a),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3a86a6),
	.w1(32'h3b8206ea),
	.w2(32'h3b23f8ba),
	.w3(32'h3aaa93ad),
	.w4(32'h3a424a61),
	.w5(32'h3b89fbfe),
	.w6(32'h3ad546ad),
	.w7(32'h3ac5f790),
	.w8(32'h3ba10fa4),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb383b7b),
	.w1(32'hbb51dcfc),
	.w2(32'hba68e852),
	.w3(32'hbb3a7615),
	.w4(32'hbb1b4b14),
	.w5(32'h364dee33),
	.w6(32'hba82d248),
	.w7(32'hbb7b14b8),
	.w8(32'h3aa73aab),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c23b251),
	.w1(32'h3bbcf423),
	.w2(32'h3ba59c22),
	.w3(32'h3c470e6e),
	.w4(32'h3bcdcca5),
	.w5(32'h3bbd15b2),
	.w6(32'h3c34185c),
	.w7(32'h3bf4aa07),
	.w8(32'h3c03b9ce),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b51b602),
	.w1(32'h3adb1c1a),
	.w2(32'h3b91e8fd),
	.w3(32'h3b93454d),
	.w4(32'h3b4b6031),
	.w5(32'h3bfeb0d8),
	.w6(32'h3bc81388),
	.w7(32'h3c0ceeec),
	.w8(32'h3b8fc2ec),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba31e386),
	.w1(32'hb8840055),
	.w2(32'h3983c72c),
	.w3(32'hbb0d2ffb),
	.w4(32'hbb0a4feb),
	.w5(32'hb804de91),
	.w6(32'hba1600e5),
	.w7(32'hbac85b8e),
	.w8(32'hba2c681f),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb06bf0d),
	.w1(32'h39ad1bb1),
	.w2(32'hba91130f),
	.w3(32'hbb09868d),
	.w4(32'h3b1dad10),
	.w5(32'h3ac2a112),
	.w6(32'hbb2a873f),
	.w7(32'hbaa02758),
	.w8(32'h3b518eca),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b104225),
	.w1(32'h3ac73501),
	.w2(32'h3b3a95b7),
	.w3(32'h399cf6dd),
	.w4(32'h3ac7e876),
	.w5(32'h3ba9738a),
	.w6(32'h3a7af5ff),
	.w7(32'h3b92ae87),
	.w8(32'h3b7b1143),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b060907),
	.w1(32'h39acca98),
	.w2(32'h3a117747),
	.w3(32'h3b443d98),
	.w4(32'h3a7b71b0),
	.w5(32'h3b3a71ac),
	.w6(32'h39265987),
	.w7(32'h3ab276b6),
	.w8(32'hbb46665f),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd5aae4),
	.w1(32'h3b4f5f66),
	.w2(32'h3c07e818),
	.w3(32'hbc0199bf),
	.w4(32'hbb5848f2),
	.w5(32'hbb162a6b),
	.w6(32'h3a8412a2),
	.w7(32'h3c107ffe),
	.w8(32'h3c7b99e6),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb884de0),
	.w1(32'h3884c5a2),
	.w2(32'h3b4769c7),
	.w3(32'hbbd2bc8e),
	.w4(32'hbba9fdc6),
	.w5(32'hb994fbe8),
	.w6(32'h3a293316),
	.w7(32'h39d361db),
	.w8(32'h3b281eef),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aee79b8),
	.w1(32'h3a3547bc),
	.w2(32'h3a7e8e6d),
	.w3(32'h3ae292ef),
	.w4(32'h3a549560),
	.w5(32'h3a978716),
	.w6(32'h3a5aec7a),
	.w7(32'h392c91a9),
	.w8(32'hba416a99),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3910d65e),
	.w1(32'hbab4d933),
	.w2(32'h39daa8b8),
	.w3(32'hbae97ebf),
	.w4(32'h397ff7dd),
	.w5(32'h3b275d3c),
	.w6(32'hbaa0d695),
	.w7(32'hbabf4471),
	.w8(32'h39e18783),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a914f7a),
	.w1(32'h3aa4435f),
	.w2(32'hb9dbc72c),
	.w3(32'hb9c7e54c),
	.w4(32'h38cc243c),
	.w5(32'hbace4be2),
	.w6(32'h3afa2f7e),
	.w7(32'hbab9b76b),
	.w8(32'hba09fd7a),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e1c245),
	.w1(32'h3894e18d),
	.w2(32'h3a319253),
	.w3(32'hbb0df8a1),
	.w4(32'h39f4c6a6),
	.w5(32'hb939e0ce),
	.w6(32'hbb3514a4),
	.w7(32'hbb33e1fb),
	.w8(32'h3ad825b6),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1f8667),
	.w1(32'hba38f0f6),
	.w2(32'h3a6e2765),
	.w3(32'h3a0ba136),
	.w4(32'hb955bc69),
	.w5(32'h3aa99416),
	.w6(32'h3b1f19d3),
	.w7(32'h3b2595d4),
	.w8(32'h3b85407c),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb288d8),
	.w1(32'hb9e668c2),
	.w2(32'h3b866fe0),
	.w3(32'h3bea15f5),
	.w4(32'h39590527),
	.w5(32'h3b7c5fd7),
	.w6(32'h3b8066de),
	.w7(32'h3b955049),
	.w8(32'h3af96826),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8b1b82),
	.w1(32'hba41cb4c),
	.w2(32'h3aabb16b),
	.w3(32'hbb2bd8ff),
	.w4(32'hbb1f3ba6),
	.w5(32'hba5f71af),
	.w6(32'hbb08580b),
	.w7(32'hbacb9cc3),
	.w8(32'hbac5ab46),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba863f42),
	.w1(32'hba850d65),
	.w2(32'hbac2fd76),
	.w3(32'hbb13cc23),
	.w4(32'hbace82b1),
	.w5(32'hbb0706f8),
	.w6(32'hbb571250),
	.w7(32'hbb16f087),
	.w8(32'hb7c34ddb),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b90ed9e),
	.w1(32'h3b04be55),
	.w2(32'h3b079041),
	.w3(32'h3badd7fb),
	.w4(32'h3b2e9411),
	.w5(32'h3affb51f),
	.w6(32'h3ba98bc3),
	.w7(32'h3b43d9bd),
	.w8(32'h3b9089b4),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9a1f6f),
	.w1(32'hba8ac599),
	.w2(32'h3aee1ec9),
	.w3(32'h3b3ca51d),
	.w4(32'hb9bd8385),
	.w5(32'hb8eb440d),
	.w6(32'h3ae1c83f),
	.w7(32'h3b110337),
	.w8(32'hbb011c2b),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9f60ed),
	.w1(32'h39e3f559),
	.w2(32'hba54927d),
	.w3(32'hbb15d98a),
	.w4(32'hba518d62),
	.w5(32'hbab3e104),
	.w6(32'hbaa2da83),
	.w7(32'hbb01783d),
	.w8(32'h3a868891),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b816dcd),
	.w1(32'h3b05344d),
	.w2(32'h3b1aea0f),
	.w3(32'h3b7d861b),
	.w4(32'h3b2f3991),
	.w5(32'h3b77fd9b),
	.w6(32'h3b95187b),
	.w7(32'h3b834bf7),
	.w8(32'h3a635a7e),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2b95f5),
	.w1(32'hbbcc3c84),
	.w2(32'hbb842eba),
	.w3(32'h39a4bac9),
	.w4(32'h3bac11ab),
	.w5(32'h3b5b6f9d),
	.w6(32'h3ba85b89),
	.w7(32'h37c17509),
	.w8(32'h39f4567e),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb0cf46),
	.w1(32'h3bacd6f3),
	.w2(32'h3cb41d2f),
	.w3(32'hbbcb745e),
	.w4(32'hbc9ec730),
	.w5(32'h3bc7d070),
	.w6(32'hbc08878d),
	.w7(32'hbc86c17b),
	.w8(32'h3b01d036),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3ae8ea),
	.w1(32'h3bb89577),
	.w2(32'h3bcb4913),
	.w3(32'h3a1eb785),
	.w4(32'h3b38252c),
	.w5(32'h3a75d0b7),
	.w6(32'h3aa7ea44),
	.w7(32'hba8fa97d),
	.w8(32'hbb0b5747),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdfde59),
	.w1(32'hbbd0f8ef),
	.w2(32'hba3e1576),
	.w3(32'hba90592f),
	.w4(32'hba1f3ec4),
	.w5(32'hb9d77e98),
	.w6(32'hbbd45207),
	.w7(32'hbbd56e22),
	.w8(32'hbb93d951),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0c4ec2),
	.w1(32'hb9de3481),
	.w2(32'hbb95d11b),
	.w3(32'hbbbb2945),
	.w4(32'h3bc06c28),
	.w5(32'h3a9be872),
	.w6(32'hba082881),
	.w7(32'hbbfb1114),
	.w8(32'hbb9af81a),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b350d9c),
	.w1(32'h3cc4cc4a),
	.w2(32'h3c670fb2),
	.w3(32'h3bf5002e),
	.w4(32'hbb22ffa2),
	.w5(32'hbbdee697),
	.w6(32'hbc231ff4),
	.w7(32'hbca1ed15),
	.w8(32'hbc065080),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1e9615),
	.w1(32'hbc4e34c6),
	.w2(32'hbc766751),
	.w3(32'hbc2a3b06),
	.w4(32'hbb94fb5e),
	.w5(32'hbbe45b04),
	.w6(32'h3a001490),
	.w7(32'hbbf69296),
	.w8(32'h3a6efe1b),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a81b708),
	.w1(32'hbb4029db),
	.w2(32'h3c042db7),
	.w3(32'h3a5716f5),
	.w4(32'hbb39ef91),
	.w5(32'h3b8194d5),
	.w6(32'hbad21f5c),
	.w7(32'h3be734c3),
	.w8(32'hba8fa234),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5639a2),
	.w1(32'hbbac5337),
	.w2(32'hbab6f569),
	.w3(32'h3ab19836),
	.w4(32'h3b73bbba),
	.w5(32'h3a510a6d),
	.w6(32'hba12426e),
	.w7(32'hbb927a6d),
	.w8(32'h3a347a39),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb9d070),
	.w1(32'h3b148a74),
	.w2(32'h3af9662d),
	.w3(32'h3be52c2e),
	.w4(32'h3ba2b0bb),
	.w5(32'h3b8b9be3),
	.w6(32'h3befe4af),
	.w7(32'h3b27df83),
	.w8(32'h3bb955ed),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c34c290),
	.w1(32'h3bfec312),
	.w2(32'h3c268af8),
	.w3(32'h3c15e39e),
	.w4(32'h3c0f5686),
	.w5(32'h3c30dcff),
	.w6(32'h3c22c19b),
	.w7(32'h3baf72fb),
	.w8(32'hba21bdd7),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9d455f),
	.w1(32'h3a80ac8d),
	.w2(32'hbb54060a),
	.w3(32'h3bba0626),
	.w4(32'hbc2eb80e),
	.w5(32'hbc09ea65),
	.w6(32'hbc8b22db),
	.w7(32'hbaa763c7),
	.w8(32'h3b3391f8),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4928b5),
	.w1(32'hb90b2e6f),
	.w2(32'hbbb67711),
	.w3(32'h3a16a9d8),
	.w4(32'h3b80606e),
	.w5(32'hba76a2ea),
	.w6(32'hba81089f),
	.w7(32'h3b055d4e),
	.w8(32'hbbebb695),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe479a1),
	.w1(32'h3bf6dbe5),
	.w2(32'hbc1b7b0a),
	.w3(32'hbc6ce56a),
	.w4(32'hbc8c8fc1),
	.w5(32'hbaee0e41),
	.w6(32'hbcd7cd7b),
	.w7(32'hbc96bfdf),
	.w8(32'hbae0dcda),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c089cfb),
	.w1(32'h3d6776a6),
	.w2(32'h3b3a4022),
	.w3(32'hbb3d4be8),
	.w4(32'h3ad617ad),
	.w5(32'h3b3099ec),
	.w6(32'h3c7ca45b),
	.w7(32'h3b205db0),
	.w8(32'hbbb64494),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b669e5d),
	.w1(32'h3d07c754),
	.w2(32'h3c12db61),
	.w3(32'hbb15577a),
	.w4(32'hbc0bcc9d),
	.w5(32'hbc8679ee),
	.w6(32'hbbffcf72),
	.w7(32'h3c20a555),
	.w8(32'h3c48c1ed),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2653c3),
	.w1(32'h3d4729d3),
	.w2(32'hbc1a43a0),
	.w3(32'hbbb1c948),
	.w4(32'hbc9afc76),
	.w5(32'h3a1de135),
	.w6(32'hbb1ac824),
	.w7(32'hbc2661e3),
	.w8(32'h3b13797f),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba52131),
	.w1(32'hba93bd27),
	.w2(32'h3c0f72f8),
	.w3(32'h3b1508b7),
	.w4(32'hbb06ef6d),
	.w5(32'h3bb6e235),
	.w6(32'hbbda879c),
	.w7(32'h3b61a9bf),
	.w8(32'hbba70cae),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2ec2b6),
	.w1(32'hbb0becc6),
	.w2(32'hbb957896),
	.w3(32'hbb53fb53),
	.w4(32'hbbcf8a56),
	.w5(32'hbc56ba8f),
	.w6(32'hbbdaa14c),
	.w7(32'hbbdd541b),
	.w8(32'h3b51b17e),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe2554a),
	.w1(32'h3c8c84d6),
	.w2(32'h3c9c3ce6),
	.w3(32'hbb495f06),
	.w4(32'h3d314f8b),
	.w5(32'h3b4ab14c),
	.w6(32'hbba9f594),
	.w7(32'h3a02e257),
	.w8(32'hbc0cfc19),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc067a27),
	.w1(32'hba513008),
	.w2(32'hbbf7e70a),
	.w3(32'hbc336afc),
	.w4(32'hba5e144a),
	.w5(32'hbc0acdbf),
	.w6(32'hbb6a9761),
	.w7(32'hbb81fd99),
	.w8(32'hbb3643a3),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe16df7),
	.w1(32'hbc0a5e3f),
	.w2(32'h39cd86d0),
	.w3(32'h3ab7bb4d),
	.w4(32'h3b62eb61),
	.w5(32'h3bb796b4),
	.w6(32'h39a74bf3),
	.w7(32'h3961997e),
	.w8(32'h3c4791d1),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c00569e),
	.w1(32'h3d0cd20e),
	.w2(32'h3c1c9333),
	.w3(32'hbb1dc8e4),
	.w4(32'hbbd11661),
	.w5(32'h3b4785ed),
	.w6(32'h3cbd4f0e),
	.w7(32'hbcbd1bb0),
	.w8(32'hba8aac89),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb37231),
	.w1(32'hbb55bab3),
	.w2(32'hbb8076c5),
	.w3(32'hbb74af04),
	.w4(32'hbb3dcc51),
	.w5(32'hbb779eb1),
	.w6(32'hb9e5705b),
	.w7(32'hbb3c3865),
	.w8(32'h3a3b023d),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b535745),
	.w1(32'h3b593884),
	.w2(32'h3aa85f6e),
	.w3(32'h3b4b75c8),
	.w4(32'h3b82ee82),
	.w5(32'h3ab003d4),
	.w6(32'h3b4d0652),
	.w7(32'h3a340875),
	.w8(32'h3ae8298d),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3958f47f),
	.w1(32'hbb3a1503),
	.w2(32'hbadea471),
	.w3(32'h3b1d52d0),
	.w4(32'h39cd5a16),
	.w5(32'hb970bd27),
	.w6(32'h3b74e7b7),
	.w7(32'h3a415ab1),
	.w8(32'h3c83a620),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c954815),
	.w1(32'hbab722e9),
	.w2(32'h3c505abd),
	.w3(32'hbba3b40e),
	.w4(32'hbc42c685),
	.w5(32'h3a32a7eb),
	.w6(32'h3c424744),
	.w7(32'h3c00c4e2),
	.w8(32'hbb02b992),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390ec233),
	.w1(32'hbb00460d),
	.w2(32'hb86341d0),
	.w3(32'h3b37f225),
	.w4(32'h3b80446e),
	.w5(32'h3ad1ad63),
	.w6(32'h39f14a00),
	.w7(32'hbac5c6c7),
	.w8(32'hbac2a295),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be16939),
	.w1(32'h3b016381),
	.w2(32'h3c2448be),
	.w3(32'hbb1d26e9),
	.w4(32'hbb8fa5e9),
	.w5(32'h3ba24584),
	.w6(32'hbc629afc),
	.w7(32'hbb928c21),
	.w8(32'h3b226107),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb31b828),
	.w1(32'hbb635a3b),
	.w2(32'hbb441ae9),
	.w3(32'h3b301849),
	.w4(32'h3b852727),
	.w5(32'h3b11ae4c),
	.w6(32'h3b20fb3d),
	.w7(32'hba86e86c),
	.w8(32'hbb4019bc),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b24a10d),
	.w1(32'hbadce5cc),
	.w2(32'h3a30ef84),
	.w3(32'h3a4bb6a5),
	.w4(32'h3b38e4bf),
	.w5(32'h3b8b8ae1),
	.w6(32'h3b6c7832),
	.w7(32'hba2a8a57),
	.w8(32'h3ba6d3c7),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e30844),
	.w1(32'hba193c17),
	.w2(32'hbae44bfc),
	.w3(32'h3b9a1298),
	.w4(32'h3b929f8a),
	.w5(32'h3ad16a63),
	.w6(32'h3b1b7aa1),
	.w7(32'hbad0337a),
	.w8(32'h3a62d4be),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ced4705),
	.w1(32'h3d3ccac3),
	.w2(32'h3c6c7f44),
	.w3(32'h3a456fb8),
	.w4(32'h3bd44293),
	.w5(32'h3c0f9bb2),
	.w6(32'h3ba63420),
	.w7(32'h3be91647),
	.w8(32'h3b064129),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab38687),
	.w1(32'hba8d329a),
	.w2(32'hbb3edf25),
	.w3(32'hbb1afa38),
	.w4(32'h3b0fb0b9),
	.w5(32'h3b8820ec),
	.w6(32'h3a04ff36),
	.w7(32'hbb6edbed),
	.w8(32'h3a90db85),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b919e19),
	.w1(32'h3b33b44a),
	.w2(32'h3bb74e2d),
	.w3(32'h3bbfb6e5),
	.w4(32'h3bb8b290),
	.w5(32'h3b9d4921),
	.w6(32'h3c03f13b),
	.w7(32'h3b5197d5),
	.w8(32'h3af12f2b),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa7d98b),
	.w1(32'hbab15842),
	.w2(32'hbb0d009b),
	.w3(32'hba559c20),
	.w4(32'h3b330f07),
	.w5(32'h3a570a56),
	.w6(32'hbaf6d117),
	.w7(32'hbb5c96b4),
	.w8(32'hbb811b64),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c17a0f9),
	.w1(32'hb8d997d7),
	.w2(32'h3c340f76),
	.w3(32'h3a3273fd),
	.w4(32'hbbacef14),
	.w5(32'h3bbb8ab9),
	.w6(32'hbc56d994),
	.w7(32'hbb9fb1ed),
	.w8(32'h3b56fa60),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbc66e0),
	.w1(32'h3b33b08b),
	.w2(32'h3bd1ec5c),
	.w3(32'h3b5f29c3),
	.w4(32'h3b121837),
	.w5(32'h3b7293a9),
	.w6(32'h3ada229d),
	.w7(32'h3ae96e1d),
	.w8(32'h3aecf4c3),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba83beae),
	.w1(32'h3ae61c6d),
	.w2(32'hbabdcd51),
	.w3(32'h399fd04a),
	.w4(32'hbb3abdca),
	.w5(32'hbb718abd),
	.w6(32'hbb6d54ff),
	.w7(32'hbb2ad9f0),
	.w8(32'hbb61271f),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c68a193),
	.w1(32'h3c14cb37),
	.w2(32'hbb71d4bb),
	.w3(32'h3ca043da),
	.w4(32'h3cbce783),
	.w5(32'h3c8e6d27),
	.w6(32'h3a2bf246),
	.w7(32'h3baaabba),
	.w8(32'hbb62b350),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4d04e3),
	.w1(32'h3b38b431),
	.w2(32'h3a8dd2af),
	.w3(32'h3b2d4d4f),
	.w4(32'h3ba32e57),
	.w5(32'h3b46601d),
	.w6(32'h3b89e316),
	.w7(32'h3a79f466),
	.w8(32'h3a35a880),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fea6d6),
	.w1(32'h3bb50d93),
	.w2(32'hbb47d360),
	.w3(32'hbac63d60),
	.w4(32'h3bc1f70c),
	.w5(32'h39aed486),
	.w6(32'hbb5bfa0c),
	.w7(32'hbbc23720),
	.w8(32'hbc9e9622),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9fa7f4),
	.w1(32'h3cdf532e),
	.w2(32'hbcc1f5a4),
	.w3(32'hbc33f344),
	.w4(32'hbc901c49),
	.w5(32'hbc02d656),
	.w6(32'hbb2154df),
	.w7(32'hbbea2c57),
	.w8(32'h3c3451a5),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b401c7f),
	.w1(32'h3bb70527),
	.w2(32'h3b3adac0),
	.w3(32'h3b595654),
	.w4(32'h3bb80c56),
	.w5(32'h3b6205e2),
	.w6(32'h3be08401),
	.w7(32'h3c0409bd),
	.w8(32'h3bb517a6),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb72f845),
	.w1(32'hbb9d5ab2),
	.w2(32'h3b4c085c),
	.w3(32'hb948abe5),
	.w4(32'h3b7e5644),
	.w5(32'h3b2e01e5),
	.w6(32'hbb2faa25),
	.w7(32'h38dcf816),
	.w8(32'h3a2a3853),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb978c549),
	.w1(32'hbb4c488a),
	.w2(32'h3c01155c),
	.w3(32'h3a661c6f),
	.w4(32'hbae60372),
	.w5(32'h3b759403),
	.w6(32'hbb84e12d),
	.w7(32'h3c20c580),
	.w8(32'hbb893a17),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a035a),
	.w1(32'hb9bbc0e2),
	.w2(32'hbb2e50b3),
	.w3(32'hbb96e5da),
	.w4(32'hbb2ecc97),
	.w5(32'hbb94017e),
	.w6(32'h38be41de),
	.w7(32'hbbaded79),
	.w8(32'hbae343c5),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaac4b0),
	.w1(32'hbbce664a),
	.w2(32'hbc1f080a),
	.w3(32'hbb6d83d1),
	.w4(32'h3ba6c501),
	.w5(32'hba8207e7),
	.w6(32'h3c38ca8f),
	.w7(32'h3a92c569),
	.w8(32'hba66b38e),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb19d5b0),
	.w1(32'hbb9362f3),
	.w2(32'h3bcea20d),
	.w3(32'hbb0ab0a2),
	.w4(32'hbb817d20),
	.w5(32'h3acebba0),
	.w6(32'hbbb1bee6),
	.w7(32'h3c00a8ef),
	.w8(32'hbb195c10),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9aa8730),
	.w1(32'hbb534ecc),
	.w2(32'h3bc5702b),
	.w3(32'h3a39af32),
	.w4(32'hbaffb28c),
	.w5(32'h3b38a669),
	.w6(32'hbb39ae3e),
	.w7(32'h3bfd37e7),
	.w8(32'h3ae92ad5),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbec6acd),
	.w1(32'hbbd9eb48),
	.w2(32'hbb837f54),
	.w3(32'hb75f940a),
	.w4(32'h3aec8016),
	.w5(32'hb9f917de),
	.w6(32'h3af5e8f7),
	.w7(32'h3b620601),
	.w8(32'hbc16eb96),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0405c8),
	.w1(32'h3b50ea99),
	.w2(32'hbc7a6551),
	.w3(32'h3c0b87a1),
	.w4(32'hbccd183f),
	.w5(32'hbc9c55ea),
	.w6(32'hbcb2fd7a),
	.w7(32'hbb22ee87),
	.w8(32'h3b2965e4),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b95ddac),
	.w1(32'h3ac1319e),
	.w2(32'h3b61c36c),
	.w3(32'h3b591fb5),
	.w4(32'h3aeb4b61),
	.w5(32'h3b816230),
	.w6(32'h3b32121a),
	.w7(32'h3a2096a4),
	.w8(32'hbac35e3a),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d299127),
	.w1(32'h3d80a6ee),
	.w2(32'h3d2d6a85),
	.w3(32'h3856b570),
	.w4(32'h3c45b929),
	.w5(32'h3c20d698),
	.w6(32'hbc7a54aa),
	.w7(32'h3c125122),
	.w8(32'h3c3fae66),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7d2d14),
	.w1(32'hbc694e54),
	.w2(32'hbc70ff89),
	.w3(32'hb9b74d79),
	.w4(32'h3bd37200),
	.w5(32'hbb32bc19),
	.w6(32'h3c5a12d4),
	.w7(32'h3c80fdec),
	.w8(32'hbbb40683),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cf84a5f),
	.w1(32'h3cd16e29),
	.w2(32'h3cf2040b),
	.w3(32'hba069138),
	.w4(32'h3c646bf0),
	.w5(32'h3c5363f9),
	.w6(32'h3c9e16a6),
	.w7(32'h3c538c5f),
	.w8(32'h3cafbf5e),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c899327),
	.w1(32'h3d4159cd),
	.w2(32'h3cad53ec),
	.w3(32'h3a756770),
	.w4(32'h3ada197b),
	.w5(32'h3be0461e),
	.w6(32'h3d85a5f9),
	.w7(32'h3cc80e06),
	.w8(32'hbb64f487),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0bcb35),
	.w1(32'hb9be2019),
	.w2(32'h3bda79fa),
	.w3(32'h3b1de31c),
	.w4(32'hbb776c6b),
	.w5(32'h3b4f0eef),
	.w6(32'hbc3e1515),
	.w7(32'hbb9d78ba),
	.w8(32'hbb10f607),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb97d14b),
	.w1(32'h39afbf4f),
	.w2(32'hba525a39),
	.w3(32'hbadb4e3b),
	.w4(32'hba971f3c),
	.w5(32'hbb5a2383),
	.w6(32'hba85183e),
	.w7(32'hbbc97608),
	.w8(32'hbbc81e06),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba021223),
	.w1(32'hbb0ba1e7),
	.w2(32'hbc6d9538),
	.w3(32'hbc04de7d),
	.w4(32'hbb2b848d),
	.w5(32'hbc965d7d),
	.w6(32'hbb9b4786),
	.w7(32'hbc35c35d),
	.w8(32'h3aee2ae3),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2ea4e7),
	.w1(32'hbb1e5b9a),
	.w2(32'hbb0d7072),
	.w3(32'h3b83938d),
	.w4(32'h3b76f216),
	.w5(32'h3b53acff),
	.w6(32'h3b90edff),
	.w7(32'h3b5f24ea),
	.w8(32'h3b9de2ef),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba9ea4d),
	.w1(32'h39e33e37),
	.w2(32'h3c0f4e7d),
	.w3(32'h3c146cc5),
	.w4(32'h3c1705ed),
	.w5(32'h3c29dc24),
	.w6(32'h3bad1cb5),
	.w7(32'h3b3d6de5),
	.w8(32'h3b766215),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba819bac),
	.w1(32'hb9c69197),
	.w2(32'hbb1f2a6b),
	.w3(32'h3b962b3d),
	.w4(32'h3bb880c4),
	.w5(32'hbaafd83f),
	.w6(32'h3c3903e0),
	.w7(32'h3c03d473),
	.w8(32'h3b0063f0),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0eee60),
	.w1(32'hba77083f),
	.w2(32'h3b7eeb02),
	.w3(32'h3a41b996),
	.w4(32'hba6c8db6),
	.w5(32'h3b048c51),
	.w6(32'hb9395232),
	.w7(32'h3b72eb54),
	.w8(32'h3aa6b1b1),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b80a882),
	.w1(32'h3b936524),
	.w2(32'h3ba02ecd),
	.w3(32'h3b0eae00),
	.w4(32'h3b3bc2c9),
	.w5(32'h3b341dc7),
	.w6(32'h3b40a555),
	.w7(32'h3b6ba7b1),
	.w8(32'h3b0c062f),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba58dae),
	.w1(32'hbb9efdf9),
	.w2(32'hbb868492),
	.w3(32'hbb8d85a7),
	.w4(32'hbb9f98ae),
	.w5(32'hbb6d0ce6),
	.w6(32'hbaf8a1af),
	.w7(32'hbb150b0b),
	.w8(32'hbb2f9788),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1c4053),
	.w1(32'hb9795509),
	.w2(32'h3a1ed9c6),
	.w3(32'h3b3c32e0),
	.w4(32'h39140afe),
	.w5(32'h3a5cd09e),
	.w6(32'h3b7db7b8),
	.w7(32'h3b0457aa),
	.w8(32'h3b00a950),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa02607),
	.w1(32'hb92ab20c),
	.w2(32'h3ac5f33d),
	.w3(32'h3ace7d3d),
	.w4(32'hba807337),
	.w5(32'h39faf189),
	.w6(32'h3b168fec),
	.w7(32'hb9669b06),
	.w8(32'h3aced0a5),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4d2eaa),
	.w1(32'h3a98406c),
	.w2(32'h3b09d523),
	.w3(32'h3b7a9d3e),
	.w4(32'h3b01b6dd),
	.w5(32'h3b3ee0d3),
	.w6(32'h3bbdf762),
	.w7(32'h3b91d0d7),
	.w8(32'h3b51dc8c),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8c3daf),
	.w1(32'h3a4f11e5),
	.w2(32'h3b3ae4f2),
	.w3(32'h3bc0395e),
	.w4(32'h3b1a44bb),
	.w5(32'h3b93f9cf),
	.w6(32'h3bd08476),
	.w7(32'h3b5aab33),
	.w8(32'h3bb3cc97),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baf6fc3),
	.w1(32'h3a79a38e),
	.w2(32'h3bb1faa1),
	.w3(32'h3be044a7),
	.w4(32'h3b0dd635),
	.w5(32'h3bd6a4c1),
	.w6(32'h3c0f8ca7),
	.w7(32'h3b887b01),
	.w8(32'h3c0883d8),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae202b7),
	.w1(32'hba039bc5),
	.w2(32'h3af98c70),
	.w3(32'h3a89841b),
	.w4(32'hbac4499d),
	.w5(32'h3a800ed6),
	.w6(32'h3b02e648),
	.w7(32'h3988704d),
	.w8(32'h3b2b5454),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb996016a),
	.w1(32'h39a7343a),
	.w2(32'hb8607a9f),
	.w3(32'hb9ed1037),
	.w4(32'h3914193e),
	.w5(32'hb9275900),
	.w6(32'hba67223f),
	.w7(32'hb99b9c7f),
	.w8(32'hba15ea1d),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9efa001),
	.w1(32'h39122b75),
	.w2(32'hb9c4cfcf),
	.w3(32'hba116d6f),
	.w4(32'h36d55a59),
	.w5(32'hb9d2d8b1),
	.w6(32'hba4d4c6e),
	.w7(32'hb975950d),
	.w8(32'hba26b486),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb65462b),
	.w1(32'hbb65a83e),
	.w2(32'hbb0d466b),
	.w3(32'hbb3e56a9),
	.w4(32'hbb4e29f5),
	.w5(32'hbb2757a2),
	.w6(32'hba78747f),
	.w7(32'hbaab6d54),
	.w8(32'hba97ae61),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b303d5b),
	.w1(32'h3a246c6b),
	.w2(32'h3b6e6ebc),
	.w3(32'h3b00390d),
	.w4(32'hb93efcbe),
	.w5(32'h3b361576),
	.w6(32'h3b8b23a8),
	.w7(32'h3acc2fff),
	.w8(32'h3b8fea6c),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1355e1),
	.w1(32'hb9e392e8),
	.w2(32'h3aa17d9d),
	.w3(32'h3a5dc365),
	.w4(32'hb97343e5),
	.w5(32'h3aa79152),
	.w6(32'h3af07d50),
	.w7(32'h3a2a8433),
	.w8(32'h3b036d80),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8192cc7),
	.w1(32'hb6076465),
	.w2(32'hb79f9f05),
	.w3(32'hb835fd00),
	.w4(32'hb6a30303),
	.w5(32'hb7cc00b9),
	.w6(32'hb897b2af),
	.w7(32'hb81a2f9b),
	.w8(32'hb859bb8b),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e9cae9),
	.w1(32'h3703019c),
	.w2(32'hb8a86e5c),
	.w3(32'hb8dce992),
	.w4(32'hb81c206c),
	.w5(32'hb8fe4f86),
	.w6(32'hb92f0133),
	.w7(32'hb89424ee),
	.w8(32'hb93b4a6f),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399793d4),
	.w1(32'h393e62d2),
	.w2(32'h3940e7c1),
	.w3(32'h39667fa1),
	.w4(32'hb90f0d22),
	.w5(32'h389722c4),
	.w6(32'h3abfa6e9),
	.w7(32'h3a3c5d41),
	.w8(32'h3a3171cd),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b301f3a),
	.w1(32'h3b29a9ac),
	.w2(32'h3b4b0916),
	.w3(32'h3b3f7060),
	.w4(32'h3b40bf8f),
	.w5(32'h3b538b97),
	.w6(32'h3b8c3dc2),
	.w7(32'h3b60632a),
	.w8(32'h3b402149),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b10a1e7),
	.w1(32'h3a997f70),
	.w2(32'h3aa4f654),
	.w3(32'h3ab19d0a),
	.w4(32'h39863259),
	.w5(32'h3a290566),
	.w6(32'h3ae33a41),
	.w7(32'h3aa54dbc),
	.w8(32'h3a761af1),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b02011c),
	.w1(32'h38f12fd5),
	.w2(32'h3b466e1b),
	.w3(32'h3b09fb20),
	.w4(32'hba1e347c),
	.w5(32'h3ad90aed),
	.w6(32'h3ae4beb2),
	.w7(32'h391f4ed8),
	.w8(32'h3b35efd4),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afe1d78),
	.w1(32'h39efc924),
	.w2(32'h3a1cbfaf),
	.w3(32'h3b283652),
	.w4(32'h3a25c1c4),
	.w5(32'h3a979f7d),
	.w6(32'h3b2dd3db),
	.w7(32'h3aa5f05e),
	.w8(32'h3af5e8e5),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394fea5e),
	.w1(32'hbadead86),
	.w2(32'hb9067796),
	.w3(32'h3a7b50c4),
	.w4(32'hbaaf83e8),
	.w5(32'h395f41eb),
	.w6(32'h3b3b46d2),
	.w7(32'h3a296f89),
	.w8(32'h3a616c8c),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37265bce),
	.w1(32'h398d0a1a),
	.w2(32'h3a410ba5),
	.w3(32'h3a342198),
	.w4(32'h39b7c411),
	.w5(32'h3ade2aaa),
	.w6(32'h3a14b0ad),
	.w7(32'h3a8edaaf),
	.w8(32'h3a98c3e2),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8bbe56),
	.w1(32'hbb0585dd),
	.w2(32'hbac235c8),
	.w3(32'hbabee661),
	.w4(32'hbaf8eb4a),
	.w5(32'hbaab51de),
	.w6(32'hba4ceaec),
	.w7(32'hbaa72207),
	.w8(32'hba344aff),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule