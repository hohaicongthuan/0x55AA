module layer_8_featuremap_221(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbad4424),
	.w1(32'h3bdaed31),
	.w2(32'h3a8885ff),
	.w3(32'hbb27659d),
	.w4(32'h3c7e262a),
	.w5(32'h3c2c52cf),
	.w6(32'h3c2cc449),
	.w7(32'h3c676aae),
	.w8(32'h3c3530ec),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aee8886),
	.w1(32'h362f521a),
	.w2(32'hbbe5edd2),
	.w3(32'h3b7df185),
	.w4(32'h3a79118b),
	.w5(32'hbb9ec76a),
	.w6(32'h3b7f69e4),
	.w7(32'hb94d16a2),
	.w8(32'h39cadf81),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf669a7),
	.w1(32'hbbb0f426),
	.w2(32'hb901ebea),
	.w3(32'hbba6b3ee),
	.w4(32'hbb952f0a),
	.w5(32'hbb9a11df),
	.w6(32'hbc40a2be),
	.w7(32'hbc2b08d4),
	.w8(32'hbb4c9f69),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b347356),
	.w1(32'h3b31b1e3),
	.w2(32'h3bebf230),
	.w3(32'h3c0eb331),
	.w4(32'h3c4f4ccf),
	.w5(32'h3c4c357d),
	.w6(32'h3b12901c),
	.w7(32'h3aee1d21),
	.w8(32'h3bec6676),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4f797b),
	.w1(32'hbcf27e36),
	.w2(32'hbd3740f8),
	.w3(32'h3b2c1aca),
	.w4(32'hbca67a8d),
	.w5(32'hbd0a5568),
	.w6(32'hbc2c5b58),
	.w7(32'hbcba2c50),
	.w8(32'hbc6c0e99),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0f48aa),
	.w1(32'h39d58c93),
	.w2(32'h3c55315e),
	.w3(32'hbcc2a911),
	.w4(32'hbac310d4),
	.w5(32'h3ae42038),
	.w6(32'hbaf97cbe),
	.w7(32'h3b8a05ca),
	.w8(32'h3a91d679),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b621077),
	.w1(32'hbc280c5c),
	.w2(32'hbbd0f5c6),
	.w3(32'h3bf0a97d),
	.w4(32'hbbd2a54b),
	.w5(32'hbb543439),
	.w6(32'hbc00ca58),
	.w7(32'hbc038be0),
	.w8(32'hbbbcf200),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb99186b),
	.w1(32'hbc065ace),
	.w2(32'hbb8ed7a5),
	.w3(32'h3aa5c9e7),
	.w4(32'hbc4ceac5),
	.w5(32'hbc03f3d0),
	.w6(32'hbbd6a21b),
	.w7(32'hbba2b6b0),
	.w8(32'hbbeecf79),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1bc6a7),
	.w1(32'hbd8cbea5),
	.w2(32'hbd9f804d),
	.w3(32'hbb2cc317),
	.w4(32'hbd811ab4),
	.w5(32'hbd952138),
	.w6(32'hbd4b2728),
	.w7(32'hbd6e2269),
	.w8(32'hbd36a450),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd745cb7),
	.w1(32'h3b139720),
	.w2(32'hbc06c263),
	.w3(32'hbd55c80b),
	.w4(32'h3c68312d),
	.w5(32'h3baf8e0d),
	.w6(32'h3afa6498),
	.w7(32'hbb862c7e),
	.w8(32'hbc3304e8),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b446c2b),
	.w1(32'hbc53ff69),
	.w2(32'hbb595e06),
	.w3(32'h3c4eb757),
	.w4(32'hbc3b11bd),
	.w5(32'hbbe667a3),
	.w6(32'hbc1cf6bf),
	.w7(32'hbbe66555),
	.w8(32'hbb6f56af),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbf9890),
	.w1(32'h3c51aa9c),
	.w2(32'h3c8f344e),
	.w3(32'hbbc4bc87),
	.w4(32'h3c9c2567),
	.w5(32'h3cd70c82),
	.w6(32'h3a939446),
	.w7(32'h3c1fca95),
	.w8(32'h3c4f7d69),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c890fa0),
	.w1(32'hbc92d5e2),
	.w2(32'hbcb75877),
	.w3(32'h3cb8d9f7),
	.w4(32'hbc47c355),
	.w5(32'hbc45c894),
	.w6(32'hbc79ac97),
	.w7(32'hbc8c1bd6),
	.w8(32'hbc853e7b),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8bda3c),
	.w1(32'h3c057ba2),
	.w2(32'h3c400606),
	.w3(32'hbc0bda6e),
	.w4(32'h3c17ddab),
	.w5(32'h3c3ab123),
	.w6(32'h3b8f91e6),
	.w7(32'h3accdcf7),
	.w8(32'hbad40886),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6fb412),
	.w1(32'hbd3bb014),
	.w2(32'hbd31a63a),
	.w3(32'h3bbf2e20),
	.w4(32'hbd2f056f),
	.w5(32'hbd2ee4a3),
	.w6(32'hbd1f28fd),
	.w7(32'hbd282582),
	.w8(32'hbd1fd013),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd2c3c3b),
	.w1(32'h3ba162d8),
	.w2(32'h3bc3aa23),
	.w3(32'hbd28f68c),
	.w4(32'h3aefb575),
	.w5(32'h3a9938aa),
	.w6(32'h3b245fa8),
	.w7(32'h3c0ebc21),
	.w8(32'h3bb32b89),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b44f4c9),
	.w1(32'hbc215db3),
	.w2(32'hbc810ea7),
	.w3(32'h3814044a),
	.w4(32'hbbc06f7c),
	.w5(32'hbc2778d8),
	.w6(32'hbb002414),
	.w7(32'hbb917df8),
	.w8(32'hbc09e69d),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2eebdc),
	.w1(32'hbb557434),
	.w2(32'hbaa9a3ea),
	.w3(32'hba13e364),
	.w4(32'hbb0943eb),
	.w5(32'h3abaeac0),
	.w6(32'hbbf230c6),
	.w7(32'hbb3326a2),
	.w8(32'h3a01c041),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c89fe59),
	.w1(32'h3c918c96),
	.w2(32'h3c5348b3),
	.w3(32'h3cb292cd),
	.w4(32'h3c8f5cb7),
	.w5(32'h3c1cfd9d),
	.w6(32'h3cccde38),
	.w7(32'h3c072873),
	.w8(32'hbc24b7b4),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2a3ee5),
	.w1(32'hbc84774b),
	.w2(32'hbc7ce0ba),
	.w3(32'h3b8bdb5c),
	.w4(32'hbc46b38b),
	.w5(32'hbc28ff21),
	.w6(32'hbc2a812e),
	.w7(32'hbc36142d),
	.w8(32'hbc6c2f15),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5fb71d),
	.w1(32'hbc69da36),
	.w2(32'hbbc8e745),
	.w3(32'hbc80028a),
	.w4(32'hbb91b488),
	.w5(32'hbba5f2b3),
	.w6(32'hbb4c833e),
	.w7(32'hbbf593eb),
	.w8(32'hbbc347e3),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc415280),
	.w1(32'hbc099e23),
	.w2(32'hbb4ec0ce),
	.w3(32'hbc2b045b),
	.w4(32'hbc0de611),
	.w5(32'hbb967270),
	.w6(32'hbba29670),
	.w7(32'hbbd6e258),
	.w8(32'hbc183c55),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c390aa1),
	.w1(32'h3ae0ed09),
	.w2(32'hbba9540c),
	.w3(32'h3c45e888),
	.w4(32'h3abaab27),
	.w5(32'hbbede3a7),
	.w6(32'h3c08511a),
	.w7(32'h3c8b800b),
	.w8(32'hbc1f3142),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeafd07),
	.w1(32'hbbaa99dd),
	.w2(32'hbb2dfb0b),
	.w3(32'hbaa94b04),
	.w4(32'hba797a0d),
	.w5(32'h3adacc94),
	.w6(32'hbb430564),
	.w7(32'h3a30f099),
	.w8(32'hba883b4e),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb239ac7),
	.w1(32'hbb64e743),
	.w2(32'hbb4c487a),
	.w3(32'h3a704f4e),
	.w4(32'hbb9151b2),
	.w5(32'hbbbc3d7b),
	.w6(32'hbbeb6709),
	.w7(32'hbc0921ec),
	.w8(32'hbc0ed80c),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a92c7dc),
	.w1(32'hbbadbad5),
	.w2(32'hbc455b3f),
	.w3(32'h3bc59e4d),
	.w4(32'hbc07edf0),
	.w5(32'hbc44eef4),
	.w6(32'h3bb847da),
	.w7(32'h3c0a3034),
	.w8(32'h3c38fd4e),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac03254),
	.w1(32'h3b8c6920),
	.w2(32'h3be4d9e4),
	.w3(32'hbb5aa6c5),
	.w4(32'hb9941e49),
	.w5(32'hbb590878),
	.w6(32'h3ae47859),
	.w7(32'h3c01bdc7),
	.w8(32'h3bcf9584),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d467eae),
	.w1(32'hbb6e1cc7),
	.w2(32'hbd03496e),
	.w3(32'h3d617ced),
	.w4(32'h3d26a208),
	.w5(32'h3c07d327),
	.w6(32'h3d33e967),
	.w7(32'h3d0b625f),
	.w8(32'hbb3b9659),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcbd493),
	.w1(32'h3ccc1520),
	.w2(32'h3c9815f0),
	.w3(32'h3c2a4c63),
	.w4(32'h3cb5d082),
	.w5(32'h3c7a82d6),
	.w6(32'h3ca68adb),
	.w7(32'h3cbc8dc0),
	.w8(32'h3baeba0e),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b20f0c4),
	.w1(32'hbc7a45bb),
	.w2(32'hbcaa0987),
	.w3(32'hbb868ced),
	.w4(32'h3a905ee2),
	.w5(32'hbb284d1f),
	.w6(32'hbbf63754),
	.w7(32'hbc38c19f),
	.w8(32'h3b9cbcca),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b019bf5),
	.w1(32'h3c091309),
	.w2(32'h3c341aaa),
	.w3(32'h3c9fc65b),
	.w4(32'h3ad50cb5),
	.w5(32'h3b531210),
	.w6(32'h3bcf38b7),
	.w7(32'h3c35aaec),
	.w8(32'h3b41693d),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c05a1b6),
	.w1(32'hbb256252),
	.w2(32'h3b17aa7e),
	.w3(32'h39f6765e),
	.w4(32'hbc6fef1a),
	.w5(32'hbbb0cf41),
	.w6(32'hbbe189e8),
	.w7(32'hbb6a3639),
	.w8(32'hbc525ce5),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc26782),
	.w1(32'h3b9b04a3),
	.w2(32'h3b82e713),
	.w3(32'hbc383fd3),
	.w4(32'h3bac0e3e),
	.w5(32'h3bee264e),
	.w6(32'h3a008025),
	.w7(32'h3a7fa7eb),
	.w8(32'hb967a346),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b51b8a8),
	.w1(32'h3bf93194),
	.w2(32'h3b3eb156),
	.w3(32'h3b8fb103),
	.w4(32'h3bf3a406),
	.w5(32'h3c2c9dcf),
	.w6(32'h3b583b1d),
	.w7(32'h3b9b454c),
	.w8(32'hbb34b726),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcf7931),
	.w1(32'hbcc4e230),
	.w2(32'hbcbb873d),
	.w3(32'h3b3cbbde),
	.w4(32'h3b4ad290),
	.w5(32'h3b8a56da),
	.w6(32'hbb88face),
	.w7(32'hbb3f8cb4),
	.w8(32'h3a5e7b0b),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1a746d),
	.w1(32'h3ad0efd8),
	.w2(32'hbc165c2c),
	.w3(32'h3c690449),
	.w4(32'h3adcc29f),
	.w5(32'hbc0c5bbd),
	.w6(32'h3b238d1b),
	.w7(32'hbb339cee),
	.w8(32'hba06829c),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa88b91),
	.w1(32'h3a6819ed),
	.w2(32'hbb84c0ed),
	.w3(32'h3a429457),
	.w4(32'h3bede576),
	.w5(32'h3b0b7198),
	.w6(32'h38b99b80),
	.w7(32'hbae7c820),
	.w8(32'hbb5d7ab6),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc26838),
	.w1(32'hbcdc52ee),
	.w2(32'hbcfcd357),
	.w3(32'hbb5dbeaa),
	.w4(32'hbc8b748a),
	.w5(32'hbcbd9710),
	.w6(32'hbc63e709),
	.w7(32'hbc9aeca6),
	.w8(32'hbc1bd0cb),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8a963a),
	.w1(32'hbb20a0c0),
	.w2(32'h3b40488e),
	.w3(32'hbc105074),
	.w4(32'hbbb52d17),
	.w5(32'hb9a3c70e),
	.w6(32'hbac8b6c4),
	.w7(32'h3b09a052),
	.w8(32'h39fd9a75),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb998ffbb),
	.w1(32'hb9bc00a1),
	.w2(32'h3aa72a63),
	.w3(32'hba252800),
	.w4(32'h3aa0b504),
	.w5(32'h3bcfb4d6),
	.w6(32'hb8f2049c),
	.w7(32'h3abd3856),
	.w8(32'h3a451182),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb07c1d),
	.w1(32'h3c5305c7),
	.w2(32'h3c83ffd9),
	.w3(32'h3cb9cb5f),
	.w4(32'h3ce38710),
	.w5(32'h3ce789ff),
	.w6(32'h3cf179a4),
	.w7(32'h3cd01e66),
	.w8(32'h3cd645b2),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8f3d86),
	.w1(32'hbc347855),
	.w2(32'h39bdb272),
	.w3(32'h3ca3bbea),
	.w4(32'hbc52b4e3),
	.w5(32'h3b00d5c3),
	.w6(32'hbc0e8b2e),
	.w7(32'hbb5b4bb1),
	.w8(32'h3b1b8b2a),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7fdf4c),
	.w1(32'hbc2d5c15),
	.w2(32'hbb614c1b),
	.w3(32'h3c66c85e),
	.w4(32'hbc473005),
	.w5(32'hbb9e62e2),
	.w6(32'hbc733c5e),
	.w7(32'hbba2903d),
	.w8(32'hbba2e916),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6ecbd5),
	.w1(32'hb9db884e),
	.w2(32'h3a8e7be4),
	.w3(32'h3ad62dd4),
	.w4(32'h3a6f8a77),
	.w5(32'h3b63e2b4),
	.w6(32'h3b073422),
	.w7(32'h3bac3304),
	.w8(32'h3aaf1151),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b37a41d),
	.w1(32'hbb2e6c18),
	.w2(32'h3b8ea593),
	.w3(32'h3b4f07e0),
	.w4(32'hb9d7642a),
	.w5(32'h3aa39d6d),
	.w6(32'h3b836d8e),
	.w7(32'h3c19a1d7),
	.w8(32'h3bf831ec),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c81a9cd),
	.w1(32'hbb95fc47),
	.w2(32'hbb5d78e6),
	.w3(32'h3c3666fe),
	.w4(32'hbb8a742c),
	.w5(32'hbb9581c2),
	.w6(32'h3a8cf7ba),
	.w7(32'hbabffba4),
	.w8(32'hbc096d7b),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a88ff),
	.w1(32'hbc4fda78),
	.w2(32'hbc94a42d),
	.w3(32'hbb1f2f73),
	.w4(32'hbc40232a),
	.w5(32'hbc805742),
	.w6(32'hbbe4cb11),
	.w7(32'hbc409dbd),
	.w8(32'hbc6c5632),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc88a4d5),
	.w1(32'hbb675bee),
	.w2(32'hb9ef9c93),
	.w3(32'hbc53414c),
	.w4(32'h3adc27ac),
	.w5(32'hbbd3911a),
	.w6(32'h3aee6c6f),
	.w7(32'hbb93ed50),
	.w8(32'hbb6d5f49),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aec5e02),
	.w1(32'hbbb66344),
	.w2(32'hbb381699),
	.w3(32'hbb3d33e2),
	.w4(32'hbadbc10f),
	.w5(32'hbb55aa17),
	.w6(32'h3a01cfaf),
	.w7(32'h3b4c716a),
	.w8(32'h3b218585),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c17a9e8),
	.w1(32'h3be34855),
	.w2(32'h3c370946),
	.w3(32'h3c1a7c91),
	.w4(32'h3c61a63e),
	.w5(32'h3c187881),
	.w6(32'h3be903f7),
	.w7(32'h3b2faba3),
	.w8(32'hb997968b),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc454825),
	.w1(32'hbba60fc9),
	.w2(32'h3c114810),
	.w3(32'hbc66015e),
	.w4(32'hbca83d1f),
	.w5(32'hbb929bd9),
	.w6(32'hbc87f739),
	.w7(32'hbbde13e0),
	.w8(32'hbca1a364),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf1860e),
	.w1(32'h3ae10e64),
	.w2(32'h39d2c195),
	.w3(32'h3c102afd),
	.w4(32'h3c4cefd7),
	.w5(32'h3bcec900),
	.w6(32'h3c70d1cf),
	.w7(32'h3bc7b7bb),
	.w8(32'h3b1446ea),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba406c8),
	.w1(32'hbc69698f),
	.w2(32'hbcacef4b),
	.w3(32'h3c407c3c),
	.w4(32'hbbe6209b),
	.w5(32'hbc49124c),
	.w6(32'hbaf209bf),
	.w7(32'hbbaffd24),
	.w8(32'hbbe05097),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc810e4d),
	.w1(32'h3a5929d6),
	.w2(32'hbb9f3df7),
	.w3(32'hbc1f46c0),
	.w4(32'h3add298d),
	.w5(32'hba07c5b8),
	.w6(32'hbbb0ee4f),
	.w7(32'hbb355f4e),
	.w8(32'h3a20969c),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b06b75e),
	.w1(32'hb9b911f8),
	.w2(32'h3c3b6ad4),
	.w3(32'h3c090431),
	.w4(32'h3afb88ef),
	.w5(32'h3bb32c08),
	.w6(32'h3ab0b0e4),
	.w7(32'h3ae49ad5),
	.w8(32'h3bae89b5),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c91eef3),
	.w1(32'h3a02eb44),
	.w2(32'hbc10649a),
	.w3(32'h3c938960),
	.w4(32'h3b6f7acb),
	.w5(32'hbba2690c),
	.w6(32'h3b572c8e),
	.w7(32'h3b1577b5),
	.w8(32'hbac2cb25),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abc5453),
	.w1(32'h3bc880e6),
	.w2(32'hbb7b79b6),
	.w3(32'hb9512053),
	.w4(32'h3c36a2f4),
	.w5(32'h3bd4d5d0),
	.w6(32'h3c0d45ec),
	.w7(32'hba01d83c),
	.w8(32'h3c04ddf0),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c00e125),
	.w1(32'hbc1dec0f),
	.w2(32'hbce11175),
	.w3(32'h3c9aaf2d),
	.w4(32'hbb69c1dd),
	.w5(32'hbcd179d4),
	.w6(32'hbb60447c),
	.w7(32'hbcad2869),
	.w8(32'hbc395458),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc24321a),
	.w1(32'h3c21b0ea),
	.w2(32'h3c3840ee),
	.w3(32'hbc53857d),
	.w4(32'h3c1bb96e),
	.w5(32'h3c5b833d),
	.w6(32'h3bbf3fce),
	.w7(32'h3c3b09f5),
	.w8(32'h3bb6a489),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c714618),
	.w1(32'h3b258d89),
	.w2(32'h3b2d8a1f),
	.w3(32'h3c841864),
	.w4(32'h3938c0bf),
	.w5(32'h3c0b854d),
	.w6(32'hbb2bfe1e),
	.w7(32'h3b9be888),
	.w8(32'h3ae07651),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2690de),
	.w1(32'hb9f8ac02),
	.w2(32'h3be9f4dd),
	.w3(32'h3ac45d8b),
	.w4(32'hbc359ff1),
	.w5(32'hbbca65ca),
	.w6(32'hba27c89a),
	.w7(32'h3bc28c6b),
	.w8(32'h3ab0dc2e),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd903e3),
	.w1(32'hbc7f57d6),
	.w2(32'hbc4d2669),
	.w3(32'hbbc232f1),
	.w4(32'hbb5f9aa4),
	.w5(32'hbc070c05),
	.w6(32'hbc15ca22),
	.w7(32'hbc2cd21e),
	.w8(32'hbc0c34cc),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd20c9f),
	.w1(32'hb9cd6e7b),
	.w2(32'h3c306655),
	.w3(32'h3b08ec85),
	.w4(32'h3be4bd52),
	.w5(32'h3c8c8748),
	.w6(32'hbb8c4424),
	.w7(32'h3b808da7),
	.w8(32'h3b3daf01),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c97ce46),
	.w1(32'h3b68b3e0),
	.w2(32'hbb389db1),
	.w3(32'h3c76fd3c),
	.w4(32'h3bffd7dd),
	.w5(32'h3b047baf),
	.w6(32'h3bb50be3),
	.w7(32'hb8aad21f),
	.w8(32'h3be02723),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3988ea),
	.w1(32'h3c8828bd),
	.w2(32'h3ca2e7e3),
	.w3(32'h3c0528d0),
	.w4(32'h3c6253de),
	.w5(32'h3c871e76),
	.w6(32'h3c192826),
	.w7(32'h3c7117c7),
	.w8(32'h3c1c5004),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c41c006),
	.w1(32'h3b71236b),
	.w2(32'h3b02b9b0),
	.w3(32'h3c0eae59),
	.w4(32'h3b40aaa4),
	.w5(32'hba06afe5),
	.w6(32'h3bc82ea4),
	.w7(32'h3b2fdc64),
	.w8(32'hbaa456a9),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad0ebcd),
	.w1(32'h3acc6a5b),
	.w2(32'h3b67a001),
	.w3(32'h3b89e86e),
	.w4(32'hb9080cbf),
	.w5(32'hbbbdc320),
	.w6(32'h3bac8b40),
	.w7(32'h3aff0c3a),
	.w8(32'h3a569de3),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba3aedb),
	.w1(32'hbb54b9ff),
	.w2(32'hbc30568c),
	.w3(32'h3c139770),
	.w4(32'hbc163380),
	.w5(32'hbc0f1068),
	.w6(32'h3bc5e43e),
	.w7(32'hbab6a286),
	.w8(32'hbbc4d8aa),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc164ee4),
	.w1(32'hba9d9bf5),
	.w2(32'h3b9a2132),
	.w3(32'hbbcae853),
	.w4(32'h3a3c9b69),
	.w5(32'h3a5d7df7),
	.w6(32'h3b333d0b),
	.w7(32'h393b2fc9),
	.w8(32'h3abeb225),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c04f7dd),
	.w1(32'h3b80a761),
	.w2(32'h3c0d652b),
	.w3(32'h3c935b1b),
	.w4(32'h3c00befb),
	.w5(32'h3c4b999e),
	.w6(32'h3c5c860e),
	.w7(32'h3c380970),
	.w8(32'h3b9a0f30),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7dfd24),
	.w1(32'hbc00f336),
	.w2(32'h3b64f822),
	.w3(32'h390e08e6),
	.w4(32'hbc178bcd),
	.w5(32'hbb1f0047),
	.w6(32'hbb45bcee),
	.w7(32'hbb45938f),
	.w8(32'h3bd2eb63),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c94c54c),
	.w1(32'h3aa4626c),
	.w2(32'h3b95f564),
	.w3(32'h3ca4e117),
	.w4(32'hbacae16f),
	.w5(32'h3b60943a),
	.w6(32'h3b6a6458),
	.w7(32'h3b2ea71d),
	.w8(32'hb89d65c7),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8614c1),
	.w1(32'h3ae15c1c),
	.w2(32'h3c03ccdf),
	.w3(32'hbae8ea4a),
	.w4(32'hbb00fbcc),
	.w5(32'hbaa2fe4c),
	.w6(32'h395885ca),
	.w7(32'hba86e3b0),
	.w8(32'h3ae6c8ff),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba89adbc),
	.w1(32'hbb077b02),
	.w2(32'hbc796ba5),
	.w3(32'h39ca85d1),
	.w4(32'h3a510608),
	.w5(32'hbc8782f7),
	.w6(32'hbb10ebbf),
	.w7(32'hbc5c7467),
	.w8(32'hbbb5fc6f),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb25da13),
	.w1(32'h3bb4d3f0),
	.w2(32'h3c165a94),
	.w3(32'hbb157d95),
	.w4(32'h3b996a5b),
	.w5(32'h3ba9754b),
	.w6(32'h3bf7e23b),
	.w7(32'h3bf1e6c5),
	.w8(32'h3b85d321),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b88214d),
	.w1(32'h3bec9683),
	.w2(32'h3c22638e),
	.w3(32'h3b90250c),
	.w4(32'h3bd2ec41),
	.w5(32'h3c3c89d1),
	.w6(32'h3b6d3941),
	.w7(32'h3c193ef2),
	.w8(32'h3ac895a8),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1176f5),
	.w1(32'hbc1965cd),
	.w2(32'hbb8bab3c),
	.w3(32'h3c174804),
	.w4(32'hbb9a612b),
	.w5(32'hbb1e6c67),
	.w6(32'hbbd8ec21),
	.w7(32'hbb93f941),
	.w8(32'hbb5d84eb),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7c9b61),
	.w1(32'hbb335253),
	.w2(32'hbbdfe248),
	.w3(32'h3bddd833),
	.w4(32'h3b753b4d),
	.w5(32'hba737096),
	.w6(32'h3bcd2cd8),
	.w7(32'h3b9b7d97),
	.w8(32'hbab320d8),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0c7c0d),
	.w1(32'h3bdb0707),
	.w2(32'hbb0e0c4f),
	.w3(32'hbbbd6e3d),
	.w4(32'hbad74d8b),
	.w5(32'hbbd99abe),
	.w6(32'hbafa6950),
	.w7(32'hbbb8b4d4),
	.w8(32'hbbc1f281),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c235dd9),
	.w1(32'hbba480c7),
	.w2(32'h3abf7b1c),
	.w3(32'h3a8942e6),
	.w4(32'hbb843df0),
	.w5(32'h3b6219bb),
	.w6(32'hbbb86eee),
	.w7(32'h3b937e14),
	.w8(32'h38ceff35),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5442dd),
	.w1(32'hbb45170e),
	.w2(32'hbb3149af),
	.w3(32'hbb0a4694),
	.w4(32'hbbc6ee89),
	.w5(32'hbbb2ba47),
	.w6(32'hbbb9ee97),
	.w7(32'hbc1e1edf),
	.w8(32'hbbde1d66),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4400f2),
	.w1(32'h3ad4b2ec),
	.w2(32'h3ba25b89),
	.w3(32'hb78c13fe),
	.w4(32'h3befcf77),
	.w5(32'h3bd63e27),
	.w6(32'hba95e2d8),
	.w7(32'h3b41aa93),
	.w8(32'hba4b2f08),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2ae457),
	.w1(32'h3bd4d500),
	.w2(32'h3b49ca49),
	.w3(32'h3c72a14b),
	.w4(32'h3bd167d6),
	.w5(32'h3b60c44e),
	.w6(32'h3c5e4995),
	.w7(32'h3c07d820),
	.w8(32'hba290345),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b19b7b4),
	.w1(32'hba273191),
	.w2(32'h3a4a9146),
	.w3(32'h3c523aed),
	.w4(32'h3ac4719f),
	.w5(32'h3c4386af),
	.w6(32'h3bfac684),
	.w7(32'hb99b252c),
	.w8(32'h3b380b82),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c743a15),
	.w1(32'h3b9a9303),
	.w2(32'h3c02fdf1),
	.w3(32'h3ce18d83),
	.w4(32'h3c86ebe2),
	.w5(32'h3c2f9aa7),
	.w6(32'h3c57b6fe),
	.w7(32'h3c9498fc),
	.w8(32'h3bc0c328),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba4f684),
	.w1(32'hbb91496d),
	.w2(32'h3bb8b23a),
	.w3(32'h3c441744),
	.w4(32'h3a9384cd),
	.w5(32'h3b21aef5),
	.w6(32'hbbd6c1a4),
	.w7(32'h3b18513e),
	.w8(32'hb9b08f5a),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeae958),
	.w1(32'h3c273fcd),
	.w2(32'h3c34e19c),
	.w3(32'hbae3dae5),
	.w4(32'h3aaf6b36),
	.w5(32'h3b71216f),
	.w6(32'h3c2555dd),
	.w7(32'h3c1048b4),
	.w8(32'h3b82c8c7),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0272ec),
	.w1(32'h3bc36c4f),
	.w2(32'h3c2dce1e),
	.w3(32'h3a962478),
	.w4(32'h3c582480),
	.w5(32'h3caecbb8),
	.w6(32'hbc14d9f1),
	.w7(32'hbb3c90f9),
	.w8(32'hbb126bed),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c421fa6),
	.w1(32'hbc0743b0),
	.w2(32'hbc0b2be9),
	.w3(32'h3c932fc8),
	.w4(32'h3b8910bf),
	.w5(32'h3bb08791),
	.w6(32'h3b9bd478),
	.w7(32'h3b7c9560),
	.w8(32'hbae27988),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0125b4),
	.w1(32'h3bf237b1),
	.w2(32'h3c539e13),
	.w3(32'h3b91e6e2),
	.w4(32'h3bc4a0ed),
	.w5(32'h3be5fd8f),
	.w6(32'h3c3fcade),
	.w7(32'h3c0bc515),
	.w8(32'h3b8c15ac),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9a3a10),
	.w1(32'hb8c5f392),
	.w2(32'h3ad0e696),
	.w3(32'h3c185030),
	.w4(32'h3a65038c),
	.w5(32'h3af8e34e),
	.w6(32'hb9b0065e),
	.w7(32'hbadfb5be),
	.w8(32'hbacb8cd4),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a6a2d),
	.w1(32'h3c0a8644),
	.w2(32'h3b41e740),
	.w3(32'hbb8e4de2),
	.w4(32'h3b697cc3),
	.w5(32'h3b9204b6),
	.w6(32'h3732fe31),
	.w7(32'h3abb206e),
	.w8(32'h3a73011d),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be75025),
	.w1(32'h3bf88757),
	.w2(32'h3b6a159c),
	.w3(32'h3c2d642a),
	.w4(32'h3c384232),
	.w5(32'h3c33fc14),
	.w6(32'h3c38630d),
	.w7(32'h3c05831f),
	.w8(32'h3bfa9774),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfa2501),
	.w1(32'h3c311e0c),
	.w2(32'h3ba3e7b6),
	.w3(32'h3c371734),
	.w4(32'h3c46fb63),
	.w5(32'h3c09125a),
	.w6(32'h3c59e39f),
	.w7(32'h3c2af775),
	.w8(32'h3bdc684c),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b89f527),
	.w1(32'hbcea8dab),
	.w2(32'hbcd1ba4a),
	.w3(32'h3bb3b156),
	.w4(32'hbc9c1e44),
	.w5(32'hbc764498),
	.w6(32'hbcc578c7),
	.w7(32'hbc4a9b45),
	.w8(32'hbbec54ad),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc49ca95),
	.w1(32'hbb186424),
	.w2(32'hbc1334f7),
	.w3(32'h3abfb321),
	.w4(32'hbb6132d4),
	.w5(32'hbc057c42),
	.w6(32'h3bbee065),
	.w7(32'hba253a4a),
	.w8(32'hbbf2f99f),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d1c3b),
	.w1(32'h3a5f487c),
	.w2(32'hbb5188d3),
	.w3(32'hb9f70ac5),
	.w4(32'hbb68fe88),
	.w5(32'hbb696c52),
	.w6(32'h3c0644a3),
	.w7(32'h3a80792e),
	.w8(32'hbb54fab1),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9a7432),
	.w1(32'h3a67bc3f),
	.w2(32'h3b259f4e),
	.w3(32'hbbaf912f),
	.w4(32'hba9cfa1a),
	.w5(32'h3c024fdc),
	.w6(32'hbafb2557),
	.w7(32'h3a9bed61),
	.w8(32'h3a5ffe62),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1677d3),
	.w1(32'h3acd23e2),
	.w2(32'h3bc9d710),
	.w3(32'h3b23c8f2),
	.w4(32'h3b7d432b),
	.w5(32'h3be571fc),
	.w6(32'h3a1959c0),
	.w7(32'h3bb75583),
	.w8(32'hb7fc3bc9),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb706c67),
	.w1(32'h3b6d4a2a),
	.w2(32'h3c020a74),
	.w3(32'hba2f9044),
	.w4(32'hba82758b),
	.w5(32'hbb2bc897),
	.w6(32'hba3229bb),
	.w7(32'h3b45bddf),
	.w8(32'h3b414f05),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbd5cad),
	.w1(32'hbb978237),
	.w2(32'hbbdd160f),
	.w3(32'hba8cdb1d),
	.w4(32'hbaadfd58),
	.w5(32'hb8b7287d),
	.w6(32'hbbbf8937),
	.w7(32'hbc385f06),
	.w8(32'hbc095713),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc115b22),
	.w1(32'hbb1709ce),
	.w2(32'hbb8abbc6),
	.w3(32'hbb63661f),
	.w4(32'hbb9aa425),
	.w5(32'hbbd8b8ed),
	.w6(32'hbbc11cf2),
	.w7(32'hbbc6c956),
	.w8(32'hbb375a2f),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb422342),
	.w1(32'h3ba002ce),
	.w2(32'h3a852310),
	.w3(32'hbb8ca3eb),
	.w4(32'h3be9b25b),
	.w5(32'h3bcf6914),
	.w6(32'h3b16844a),
	.w7(32'h3b89c2c7),
	.w8(32'hbb5773b0),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b15d56f),
	.w1(32'h3c237eda),
	.w2(32'h3c11cb95),
	.w3(32'h3a9633a5),
	.w4(32'h3bc6c7b2),
	.w5(32'h3c235f13),
	.w6(32'h3b9ee745),
	.w7(32'h3bc18e28),
	.w8(32'h3a3f7034),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c337657),
	.w1(32'hbb94b558),
	.w2(32'h3adba2c9),
	.w3(32'h3c71df51),
	.w4(32'hbb59885c),
	.w5(32'h3a9c810f),
	.w6(32'h3b751025),
	.w7(32'h3b7d541a),
	.w8(32'hba92d716),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a163c72),
	.w1(32'hbc3a126d),
	.w2(32'hbb98de58),
	.w3(32'h3c2b9617),
	.w4(32'hbc0dca47),
	.w5(32'hbb2d4249),
	.w6(32'hbbe3f7e1),
	.w7(32'h3a074bb7),
	.w8(32'hbc43d494),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0fb2c9),
	.w1(32'h3bd5507c),
	.w2(32'h3bf5bbbf),
	.w3(32'hbc34e3a5),
	.w4(32'hba9c4506),
	.w5(32'h3b13a642),
	.w6(32'h3c1c70a8),
	.w7(32'h3c2a98db),
	.w8(32'h3b06e153),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2027df),
	.w1(32'hbc0b6620),
	.w2(32'hbbe0d564),
	.w3(32'hbb6c8fbe),
	.w4(32'hbbb6f7fb),
	.w5(32'hbbd2e60e),
	.w6(32'hbb40852a),
	.w7(32'hbae980d0),
	.w8(32'hb8f6689d),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb973549),
	.w1(32'hbb6bb6dc),
	.w2(32'hba0c834d),
	.w3(32'hbc031b7f),
	.w4(32'hba5ed2a8),
	.w5(32'h3a26ebd9),
	.w6(32'hbbac0910),
	.w7(32'hbba408e6),
	.w8(32'hbb0ac39e),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3accd26b),
	.w1(32'h3bbbc33f),
	.w2(32'h3b662692),
	.w3(32'h3aa34950),
	.w4(32'h3bdafe82),
	.w5(32'h3ba935a4),
	.w6(32'h3bc051cb),
	.w7(32'h3c056fa2),
	.w8(32'h3b9c8a3a),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbfcc25),
	.w1(32'hbb83605c),
	.w2(32'hbb99d5df),
	.w3(32'h3c134e95),
	.w4(32'h3b4810cb),
	.w5(32'hbbd34b62),
	.w6(32'hbaa01ab8),
	.w7(32'hbbb70bbc),
	.w8(32'hbb61cfe1),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb90760),
	.w1(32'h3cdf6d64),
	.w2(32'h3d031026),
	.w3(32'hbac2fc92),
	.w4(32'h3cd6bd45),
	.w5(32'h3cfd1cdb),
	.w6(32'h3cc58132),
	.w7(32'h3cd488cf),
	.w8(32'h3c9e82ec),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce101ec),
	.w1(32'hbc0df91d),
	.w2(32'hbbc45574),
	.w3(32'h3cd1ff4d),
	.w4(32'hbb93a8bb),
	.w5(32'h3b17ab2d),
	.w6(32'hbc2578ad),
	.w7(32'hbb868c87),
	.w8(32'hbb938ae3),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe8a167),
	.w1(32'hbbf67da4),
	.w2(32'hbc23ffd1),
	.w3(32'hbb83ef7b),
	.w4(32'hbc504133),
	.w5(32'hbc0ca68b),
	.w6(32'h3b29ef3c),
	.w7(32'h3b869434),
	.w8(32'h3addac44),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbda9fd4),
	.w1(32'hbc0f6625),
	.w2(32'hbba0c094),
	.w3(32'hbbffd481),
	.w4(32'hbb94df4c),
	.w5(32'hbaaf69e6),
	.w6(32'hbc2a6d65),
	.w7(32'hbbe75ecd),
	.w8(32'hbc055490),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb1bebf),
	.w1(32'h3c17ee36),
	.w2(32'h3c00738b),
	.w3(32'hbb365fee),
	.w4(32'h3c1ca655),
	.w5(32'h3c13aed2),
	.w6(32'h3bf7c4d9),
	.w7(32'h3c10f3de),
	.w8(32'h3bb96465),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b36938d),
	.w1(32'h3ada12d2),
	.w2(32'h3c3552a6),
	.w3(32'h3ba025b3),
	.w4(32'hbc099256),
	.w5(32'hbaa6c90d),
	.w6(32'h3b7dbea9),
	.w7(32'h3c222960),
	.w8(32'h3a8e5aae),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b085c8c),
	.w1(32'hbbb47e7e),
	.w2(32'hb9a2724e),
	.w3(32'hb8d755c8),
	.w4(32'hbb55875f),
	.w5(32'hba751489),
	.w6(32'h3b2279ef),
	.w7(32'h3b2183a1),
	.w8(32'h3a0ad8a2),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf5955c),
	.w1(32'h3aa27c52),
	.w2(32'h3bff1a69),
	.w3(32'hbb00d894),
	.w4(32'h3b455697),
	.w5(32'h3baee6ac),
	.w6(32'h3b10e1eb),
	.w7(32'h3ba9fffe),
	.w8(32'h3bb0afad),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c298b88),
	.w1(32'h3bb0a9de),
	.w2(32'hbb2e6c4e),
	.w3(32'h3b0a85d9),
	.w4(32'h3a7d0e9c),
	.w5(32'hbba70c8e),
	.w6(32'h3c0db09d),
	.w7(32'h3aaeb693),
	.w8(32'h3aab7dbe),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1cacda),
	.w1(32'hbc0c8da5),
	.w2(32'hbc3684ca),
	.w3(32'h3b5cc647),
	.w4(32'h39936b11),
	.w5(32'h3b0aca37),
	.w6(32'hbbdee378),
	.w7(32'hba9d12f4),
	.w8(32'h3af43cbe),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bdd25e),
	.w1(32'hbb8785c4),
	.w2(32'h3aafd987),
	.w3(32'hbae3f298),
	.w4(32'hbb8bb5a3),
	.w5(32'hbb5792e7),
	.w6(32'hbadfebb8),
	.w7(32'h3b2029a9),
	.w8(32'hbbfb0f08),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc34c3d2),
	.w1(32'hbc99e713),
	.w2(32'hbce2a2e4),
	.w3(32'hbc461588),
	.w4(32'hbc8f1243),
	.w5(32'hbccb38d8),
	.w6(32'hbc70cbdc),
	.w7(32'hbca2d0ad),
	.w8(32'hbc8e8a2c),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf1e69d),
	.w1(32'hbc2359ed),
	.w2(32'hbbab72b6),
	.w3(32'hbcd36ad9),
	.w4(32'hbc284498),
	.w5(32'hbb37cd9d),
	.w6(32'hbbb56c06),
	.w7(32'hbb0d4675),
	.w8(32'hbb598820),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb204994),
	.w1(32'h3b9f2de8),
	.w2(32'h3b4cf41b),
	.w3(32'hbbc34fb8),
	.w4(32'hbbedb3dd),
	.w5(32'hbbacdfa6),
	.w6(32'hbb311ab9),
	.w7(32'h3945ba37),
	.w8(32'h3bb56e3c),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb32fb8),
	.w1(32'hbb557a78),
	.w2(32'h3981c6ca),
	.w3(32'h3b5c8dab),
	.w4(32'hbbabb4f0),
	.w5(32'hbba981dc),
	.w6(32'hbbbda970),
	.w7(32'hbbdb4ae7),
	.w8(32'hbba82f35),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa7dc2f),
	.w1(32'hbafae217),
	.w2(32'hbb841265),
	.w3(32'h3a5d25d3),
	.w4(32'hbae307d3),
	.w5(32'hbb65f920),
	.w6(32'h3a5ca593),
	.w7(32'hbada1f76),
	.w8(32'hbaf9ab7b),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba775496),
	.w1(32'h3bb0ed4d),
	.w2(32'h39f896df),
	.w3(32'h3966facd),
	.w4(32'h3c251f19),
	.w5(32'h3c1ce44f),
	.w6(32'h3c1eb0e1),
	.w7(32'h3b6744d7),
	.w8(32'h3af558dc),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule