module layer_8_featuremap_209(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beb4bce),
	.w1(32'h3c5eae99),
	.w2(32'h3c160981),
	.w3(32'hbb234c59),
	.w4(32'h3b435d75),
	.w5(32'h3ac7e3ac),
	.w6(32'hb7c5d31e),
	.w7(32'h3c5b3131),
	.w8(32'h3cba5935),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1036f1),
	.w1(32'h3aad7fbe),
	.w2(32'h3b4e9196),
	.w3(32'hbc2a6e0c),
	.w4(32'h3b1b7e70),
	.w5(32'h3b829f95),
	.w6(32'h3a8948a6),
	.w7(32'hb9507497),
	.w8(32'h3a7f295b),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b56c33d),
	.w1(32'h3cd98198),
	.w2(32'h3ccee49c),
	.w3(32'h3b2061e6),
	.w4(32'h3ce2f504),
	.w5(32'h3ca2d348),
	.w6(32'h3c1bc94c),
	.w7(32'h3c329360),
	.w8(32'h3bf28864),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c702fc8),
	.w1(32'h3cad67ca),
	.w2(32'h3cb92c94),
	.w3(32'h3c3a0200),
	.w4(32'h3c6d3b35),
	.w5(32'h3ba84b8d),
	.w6(32'h3c112370),
	.w7(32'h3c1ee6c3),
	.w8(32'h3bed9c91),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be96977),
	.w1(32'hbb3538b0),
	.w2(32'hbc125717),
	.w3(32'hbbc11b05),
	.w4(32'hba8e74c2),
	.w5(32'hbb72f832),
	.w6(32'h3ae6dfcb),
	.w7(32'hbb1b4463),
	.w8(32'h3a43dc5e),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbabee6b),
	.w1(32'h3acf5eee),
	.w2(32'h3c9952c7),
	.w3(32'hbb912ac5),
	.w4(32'hbb33a70a),
	.w5(32'h3c4e8e6b),
	.w6(32'hb96a5f06),
	.w7(32'h3bb6f441),
	.w8(32'h3be14be8),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca54f55),
	.w1(32'hbb7b4879),
	.w2(32'hbc1d9d54),
	.w3(32'h3a981781),
	.w4(32'hbba67e34),
	.w5(32'hbc2c9542),
	.w6(32'hbb5c55d3),
	.w7(32'hbc04d1a5),
	.w8(32'hbbe3e769),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc00f8a3),
	.w1(32'hbc6f90e2),
	.w2(32'h3aba890a),
	.w3(32'hbc236767),
	.w4(32'hbbf37b44),
	.w5(32'hbcc04799),
	.w6(32'hbc816ad7),
	.w7(32'h3c278b4f),
	.w8(32'h3c02d358),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c324b31),
	.w1(32'h3c0dad81),
	.w2(32'h3c4c3f46),
	.w3(32'hbc5ef4bb),
	.w4(32'h3c02c36b),
	.w5(32'h3c4905be),
	.w6(32'hbbb5299f),
	.w7(32'hbbb2e950),
	.w8(32'hbbbb513a),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1ca8fb),
	.w1(32'h3c69ffeb),
	.w2(32'h3c313102),
	.w3(32'h3bbee784),
	.w4(32'h3c25e69c),
	.w5(32'h3ca83767),
	.w6(32'h3be23f11),
	.w7(32'hbbdd2c43),
	.w8(32'hbc95c7ca),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc68a81),
	.w1(32'hbc3d2a99),
	.w2(32'hbb8b0afb),
	.w3(32'h3c78dad8),
	.w4(32'hbc840ba1),
	.w5(32'hbc8f2c80),
	.w6(32'hbc5dbe00),
	.w7(32'hbbf7f935),
	.w8(32'hbb149b5a),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b71b1b3),
	.w1(32'hbc54100c),
	.w2(32'hbc82a5a1),
	.w3(32'hbc4fbbab),
	.w4(32'hbbd2d6a9),
	.w5(32'hbc9269fc),
	.w6(32'hbbaba95a),
	.w7(32'hbb87d190),
	.w8(32'h3c12c1bf),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb828079),
	.w1(32'h3c236c86),
	.w2(32'h3d05f2a2),
	.w3(32'h393cf892),
	.w4(32'h3bff0660),
	.w5(32'h3d1e1d79),
	.w6(32'hbbaacfb6),
	.w7(32'h3c251863),
	.w8(32'hbb1eacd1),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cf3f357),
	.w1(32'h3b896a7b),
	.w2(32'hbc5ec5da),
	.w3(32'h3cc55b69),
	.w4(32'h3c007a07),
	.w5(32'hbc4f194a),
	.w6(32'h3ba9ec00),
	.w7(32'hbbcb8e19),
	.w8(32'hbc4ffc02),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6b24da),
	.w1(32'hb9fbea6a),
	.w2(32'hba9e4538),
	.w3(32'hbca197d4),
	.w4(32'hba185f63),
	.w5(32'hbb0c1ac4),
	.w6(32'hbbc04b7d),
	.w7(32'hbbaa24f9),
	.w8(32'hbbb25666),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3993cccc),
	.w1(32'h3ca7bcae),
	.w2(32'h3c8d8cc2),
	.w3(32'hb9dabcff),
	.w4(32'h3c635fae),
	.w5(32'h3c8fd641),
	.w6(32'h3bbeed25),
	.w7(32'h3ba5f154),
	.w8(32'h3c45d0df),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abd1bf6),
	.w1(32'h3a664e3f),
	.w2(32'h3c440967),
	.w3(32'hbb04c8b9),
	.w4(32'h3a885c8e),
	.w5(32'h3b794d45),
	.w6(32'hbb2c6a82),
	.w7(32'h3a8b5bba),
	.w8(32'h3c10b5c6),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2c13b2),
	.w1(32'h3c1eb632),
	.w2(32'h3c42815a),
	.w3(32'h3b6b7bdb),
	.w4(32'h3c16cf6d),
	.w5(32'h3c06c2af),
	.w6(32'hbb8daf43),
	.w7(32'h3b430cf2),
	.w8(32'hbbc9f5e5),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc95814),
	.w1(32'hbc96a34c),
	.w2(32'hbcf69d2b),
	.w3(32'h3accc4a6),
	.w4(32'hbc60737b),
	.w5(32'hbccade2b),
	.w6(32'hbc522e81),
	.w7(32'hbc7a1018),
	.w8(32'hbc0ff632),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7036d6),
	.w1(32'h3be9acbd),
	.w2(32'h3c2969ab),
	.w3(32'hbc7408b6),
	.w4(32'h3bab860b),
	.w5(32'h3bd73c0a),
	.w6(32'hbb987fd7),
	.w7(32'hbb355bf0),
	.w8(32'hbbb0a6de),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbaaff1),
	.w1(32'h3c1c009c),
	.w2(32'h3c8a71dd),
	.w3(32'h3b89dbbf),
	.w4(32'h3c5961fd),
	.w5(32'h3c94a60d),
	.w6(32'h3afd7597),
	.w7(32'h3b9ab04e),
	.w8(32'hba66f705),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0504ad),
	.w1(32'h3cb54ac3),
	.w2(32'h3d27fd5a),
	.w3(32'h3bbc8890),
	.w4(32'h3cb7025d),
	.w5(32'h3cec06c7),
	.w6(32'h3c042d9d),
	.w7(32'h3cd09d33),
	.w8(32'h3c818938),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d0de3dc),
	.w1(32'h3c77d81a),
	.w2(32'h3c6857ac),
	.w3(32'h3ca230e6),
	.w4(32'h3c11ff8e),
	.w5(32'h3c4971c2),
	.w6(32'h3bb6b538),
	.w7(32'h3c3e8efb),
	.w8(32'hbb231c55),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac4c5d0),
	.w1(32'h3c8f0427),
	.w2(32'h3d0f2689),
	.w3(32'h3ba6ed9d),
	.w4(32'h3c8c8f34),
	.w5(32'h3cd7f077),
	.w6(32'h3bc68256),
	.w7(32'h3c580cdb),
	.w8(32'h3c5ddfa9),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce47d6e),
	.w1(32'h3b9c0fff),
	.w2(32'h3bf0e597),
	.w3(32'h3c5ee9fb),
	.w4(32'h3c158bf7),
	.w5(32'h3c5d6b3d),
	.w6(32'h3a1f13af),
	.w7(32'h3b4c956c),
	.w8(32'hbba65349),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac998ef),
	.w1(32'h3c404e46),
	.w2(32'h3c5ae3d9),
	.w3(32'h3ab6afdb),
	.w4(32'h3b81b553),
	.w5(32'h3af34917),
	.w6(32'h3b1b6e38),
	.w7(32'h3bd3d2ca),
	.w8(32'h3b0947f6),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba362bb),
	.w1(32'h3c9bdd0d),
	.w2(32'h3ca970e1),
	.w3(32'hba55c2c2),
	.w4(32'h3c89424e),
	.w5(32'h3c113d82),
	.w6(32'h3ae9cd90),
	.w7(32'h3ca5376a),
	.w8(32'h3c976654),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8a9c34),
	.w1(32'h3b79b08c),
	.w2(32'h3bec7314),
	.w3(32'hbbb66456),
	.w4(32'hba3d113c),
	.w5(32'h3b423d4b),
	.w6(32'hbacda1f9),
	.w7(32'hbb4fae84),
	.w8(32'hbbaae3b7),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbe27d8),
	.w1(32'hbbf657c6),
	.w2(32'hbbe3d8e4),
	.w3(32'h38476568),
	.w4(32'hbbba9939),
	.w5(32'hbb556cdc),
	.w6(32'hbc4c0d95),
	.w7(32'hbc8edb17),
	.w8(32'hbc03cb02),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a54d0ff),
	.w1(32'hbbfb9001),
	.w2(32'hbbcf705e),
	.w3(32'h3ba74d85),
	.w4(32'h3bbe4db4),
	.w5(32'hba2fbff0),
	.w6(32'hbb8978dc),
	.w7(32'hbba03d5b),
	.w8(32'h3c338778),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbeff30),
	.w1(32'h3b902e87),
	.w2(32'h3b376a34),
	.w3(32'h3c383bfb),
	.w4(32'h3bbb6f24),
	.w5(32'h3c0dcfff),
	.w6(32'h3a1f5af9),
	.w7(32'h3b10c73d),
	.w8(32'hbb4fe0be),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae088ac),
	.w1(32'h3b58d68a),
	.w2(32'h3b2c49bb),
	.w3(32'h3b92da53),
	.w4(32'h3b0c1659),
	.w5(32'h3a236b24),
	.w6(32'hbb3b1446),
	.w7(32'hbb42aa76),
	.w8(32'hbb941abb),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9a1c83),
	.w1(32'h3c33f1e9),
	.w2(32'h3c9f9ee4),
	.w3(32'h3ac55da1),
	.w4(32'h3bf1f5f9),
	.w5(32'h3b8caf77),
	.w6(32'h3bef074e),
	.w7(32'h3c06e782),
	.w8(32'hba9236ce),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baf4386),
	.w1(32'hbbac91c1),
	.w2(32'hbccada3d),
	.w3(32'h3bac06a7),
	.w4(32'hbc199dc5),
	.w5(32'hbc2e56cb),
	.w6(32'h3b621fbe),
	.w7(32'hbb553721),
	.w8(32'h3b234ff3),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3f1c29),
	.w1(32'h3acd90b0),
	.w2(32'h3bd41757),
	.w3(32'hbc46629f),
	.w4(32'hbb85fc1c),
	.w5(32'h3b909d61),
	.w6(32'hba8e15ce),
	.w7(32'hba792a57),
	.w8(32'h3c0ab0d7),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6a42d9),
	.w1(32'hbcc30f87),
	.w2(32'hbd8918d9),
	.w3(32'h3c193735),
	.w4(32'hbd262298),
	.w5(32'hbd98de59),
	.w6(32'hbc3773f8),
	.w7(32'hbca3bd4d),
	.w8(32'hbcb544fa),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd530269),
	.w1(32'h3b5ab6ea),
	.w2(32'h3c0e8cfb),
	.w3(32'hbd3b6fba),
	.w4(32'h3bacb4d1),
	.w5(32'h3c273eb8),
	.w6(32'hbb1de6e4),
	.w7(32'hb81c16c9),
	.w8(32'hb93d8104),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0039ee),
	.w1(32'h3b0b476f),
	.w2(32'h3bdaaf98),
	.w3(32'h3c47fe59),
	.w4(32'h3b0894a2),
	.w5(32'h3b8514e8),
	.w6(32'hbb4ea99e),
	.w7(32'h39e7ac4d),
	.w8(32'hbb3f7fd3),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b91ca53),
	.w1(32'h3bf1ae2c),
	.w2(32'h3bc4adc8),
	.w3(32'h3b38f8b6),
	.w4(32'h3c0adeef),
	.w5(32'h3bc0a2a7),
	.w6(32'hbb5cb853),
	.w7(32'hbc02f2b2),
	.w8(32'hbb717cfb),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c26e53e),
	.w1(32'hb9016abe),
	.w2(32'hbc052c15),
	.w3(32'h3c2ccc28),
	.w4(32'hbbc36664),
	.w5(32'hbb416173),
	.w6(32'h3b2b66b5),
	.w7(32'hb97319b7),
	.w8(32'h3b294a6c),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2fcea9),
	.w1(32'h3c0112fb),
	.w2(32'h3c6fdc81),
	.w3(32'h3b09322c),
	.w4(32'h3c0154f5),
	.w5(32'h3c633f07),
	.w6(32'h3b916cb5),
	.w7(32'h3c3b9fff),
	.w8(32'h3be223e6),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c22d455),
	.w1(32'h3bf432af),
	.w2(32'h3b97176e),
	.w3(32'h3c0df6c2),
	.w4(32'h3b96caf5),
	.w5(32'h3be4613e),
	.w6(32'hbb94850e),
	.w7(32'hbc0659c3),
	.w8(32'hbc42c9e4),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb305cf1),
	.w1(32'hbc184ccb),
	.w2(32'hbbd11910),
	.w3(32'h3b97c498),
	.w4(32'hbc09adf0),
	.w5(32'hbbae9da5),
	.w6(32'hbbd83e41),
	.w7(32'hbc02e6f9),
	.w8(32'hbc410384),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf777e7),
	.w1(32'h3a252310),
	.w2(32'h3c448bb3),
	.w3(32'hbb5cb61e),
	.w4(32'h3abffae7),
	.w5(32'h3bd2b426),
	.w6(32'hbc21a1ff),
	.w7(32'h3ba0c373),
	.w8(32'hbb5999d4),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4af290),
	.w1(32'h3b7eb362),
	.w2(32'hbc95ee03),
	.w3(32'h3c304c8f),
	.w4(32'h3b891d13),
	.w5(32'hbb9d5c1c),
	.w6(32'h3b8d22d2),
	.w7(32'hbbe90087),
	.w8(32'hbb1e1174),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc871929),
	.w1(32'h3c200b2e),
	.w2(32'h3afe4ad2),
	.w3(32'h3b5bd108),
	.w4(32'h3b9de20d),
	.w5(32'hbba0914c),
	.w6(32'h3b4ddd60),
	.w7(32'hbbbad6c9),
	.w8(32'hbb68d176),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b60a597),
	.w1(32'hbc17b5ed),
	.w2(32'hbc735ce1),
	.w3(32'hbb8fb654),
	.w4(32'hbbd56f46),
	.w5(32'hbc726016),
	.w6(32'hbbfa6996),
	.w7(32'hbc0c606f),
	.w8(32'h3a7c2b91),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcebf2d),
	.w1(32'hbc0f002c),
	.w2(32'hbd14397b),
	.w3(32'hbc3977e4),
	.w4(32'hbc38e8c2),
	.w5(32'hbd072dd1),
	.w6(32'hbba87bc2),
	.w7(32'hbc783399),
	.w8(32'hbc0691a4),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce85687),
	.w1(32'h3bf2ea44),
	.w2(32'hbc889886),
	.w3(32'hbcbb422d),
	.w4(32'h3ba04ace),
	.w5(32'hbbcf62a1),
	.w6(32'h3b037c3c),
	.w7(32'hbb89f7e7),
	.w8(32'hbbf1b1f9),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc819b07),
	.w1(32'hbbea269e),
	.w2(32'hbba1c17c),
	.w3(32'hbc111d19),
	.w4(32'h3aab3a4d),
	.w5(32'h3b3cd332),
	.w6(32'hbbd1093d),
	.w7(32'hbc450ff1),
	.w8(32'hbc3f76b6),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc806514),
	.w1(32'h3ba0f550),
	.w2(32'hbc214dc7),
	.w3(32'hbbe01248),
	.w4(32'h39dff957),
	.w5(32'hbc12e00a),
	.w6(32'h3b54e9a9),
	.w7(32'hbbace76e),
	.w8(32'h3b7ae6e4),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a06d62e),
	.w1(32'hbc0f3067),
	.w2(32'hbc1a62c8),
	.w3(32'hba225101),
	.w4(32'hbc0e7e29),
	.w5(32'hbc1738e6),
	.w6(32'hbbdfc4a4),
	.w7(32'hbc17b818),
	.w8(32'hbba5739a),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb195349),
	.w1(32'h3b3dafe2),
	.w2(32'hbb742dbc),
	.w3(32'hbbe8a065),
	.w4(32'hbb740229),
	.w5(32'hbbd87e2a),
	.w6(32'h3b902d8e),
	.w7(32'h38a131f4),
	.w8(32'h39f0de83),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadc293e),
	.w1(32'hbcd9cc06),
	.w2(32'hbc896dc1),
	.w3(32'hbc06f10b),
	.w4(32'hbc83d3bc),
	.w5(32'hbc362190),
	.w6(32'hbc8dadff),
	.w7(32'hbc3777d8),
	.w8(32'hbc022764),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1ed467),
	.w1(32'hbc33fad7),
	.w2(32'hbb0e1544),
	.w3(32'h3c2bc90c),
	.w4(32'hbc4faf78),
	.w5(32'h3891f048),
	.w6(32'h3ac52baf),
	.w7(32'h3903ae27),
	.w8(32'hbc159e9c),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2303ec),
	.w1(32'h3cc0c76b),
	.w2(32'h3d2b68fc),
	.w3(32'hbbf2ec1d),
	.w4(32'h3c752e4c),
	.w5(32'h3cdfe805),
	.w6(32'h3c00b2cf),
	.w7(32'h3cb35177),
	.w8(32'h3c7b2bdc),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cf67719),
	.w1(32'h3aaa603f),
	.w2(32'hb989c945),
	.w3(32'h3c8d3472),
	.w4(32'hbbcf02ed),
	.w5(32'hbbbb5f7e),
	.w6(32'hbb7ac593),
	.w7(32'h3ab6fef6),
	.w8(32'h3b97b1a9),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ada912e),
	.w1(32'hbbae9414),
	.w2(32'hbc106772),
	.w3(32'hb9c2d4bb),
	.w4(32'h39c54f7c),
	.w5(32'hbbce258b),
	.w6(32'hbabb74fa),
	.w7(32'hbc008574),
	.w8(32'h39692106),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b743ab2),
	.w1(32'h3b9f682b),
	.w2(32'h3ba44e63),
	.w3(32'h3bf7e659),
	.w4(32'h3be7ac59),
	.w5(32'h3b9d985a),
	.w6(32'h3b83a2ad),
	.w7(32'h3bca42cc),
	.w8(32'h3bfaa416),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb65676),
	.w1(32'h3ca85ab8),
	.w2(32'h3cf00998),
	.w3(32'h3b5c36c6),
	.w4(32'h3c72409a),
	.w5(32'h3c9c26bf),
	.w6(32'h3baba297),
	.w7(32'h3c699e1c),
	.w8(32'h3c5a7887),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cdb7348),
	.w1(32'h3c2f0a3c),
	.w2(32'h3d16ddb2),
	.w3(32'h3ca9d50e),
	.w4(32'h3c029e18),
	.w5(32'h3cea14a0),
	.w6(32'hba2cfb04),
	.w7(32'h3c355c3b),
	.w8(32'hbb1e6554),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ccae915),
	.w1(32'h3b344665),
	.w2(32'hba6f867d),
	.w3(32'h3c69eae7),
	.w4(32'h3b99e100),
	.w5(32'h3b1e9f9b),
	.w6(32'hbbb066c1),
	.w7(32'hbb779da4),
	.w8(32'hbc422545),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbb8713),
	.w1(32'h3c46f3ec),
	.w2(32'hbb3911e9),
	.w3(32'h3b0d0c33),
	.w4(32'h3bb5db1f),
	.w5(32'hbc28f69e),
	.w6(32'h3a213416),
	.w7(32'hbc4f5c7d),
	.w8(32'hbc047218),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9779af),
	.w1(32'h3b465c64),
	.w2(32'h3a94d2a6),
	.w3(32'hba4247c6),
	.w4(32'h3b481da8),
	.w5(32'h3aeed86e),
	.w6(32'h3b9f948b),
	.w7(32'h3acf34d0),
	.w8(32'hbab13918),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba93a791),
	.w1(32'h3a7437cf),
	.w2(32'h3aa5a58b),
	.w3(32'hbb7177e7),
	.w4(32'h3aaa191a),
	.w5(32'h3b372b01),
	.w6(32'h3a839215),
	.w7(32'hba3c58df),
	.w8(32'h381da5c4),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b15ad6e),
	.w1(32'h3a84c3f1),
	.w2(32'hbb888906),
	.w3(32'h3be721e0),
	.w4(32'hbb496b5f),
	.w5(32'hbc087fa4),
	.w6(32'h3b0f0431),
	.w7(32'hbc31b6c7),
	.w8(32'hbb5d791d),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafe9c36),
	.w1(32'h3b9fe79b),
	.w2(32'h3ca2ca25),
	.w3(32'hbbdbc644),
	.w4(32'h3aeaabe7),
	.w5(32'h3c8de8f7),
	.w6(32'hbac98262),
	.w7(32'h3c5ab64e),
	.w8(32'h3b3de970),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9af0e5),
	.w1(32'h3bbe2d00),
	.w2(32'h3bb82aa3),
	.w3(32'h3c4858b9),
	.w4(32'h3c3d8adf),
	.w5(32'h3bc728dc),
	.w6(32'hbbac0737),
	.w7(32'h3c25244b),
	.w8(32'h3bf922e6),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb59ab0c),
	.w1(32'h3c8e78db),
	.w2(32'h3cd18b61),
	.w3(32'h3bab65c3),
	.w4(32'h3c0d1aea),
	.w5(32'h3c6f1656),
	.w6(32'h3c3045dc),
	.w7(32'h3c540e52),
	.w8(32'h3b9f20b8),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd15edd),
	.w1(32'h3c6fb056),
	.w2(32'h3ceb5160),
	.w3(32'h3ae13815),
	.w4(32'h3c80cab2),
	.w5(32'h3cb47d62),
	.w6(32'h3aadf87d),
	.w7(32'h3bb9bde0),
	.w8(32'h3c004ce1),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c776a36),
	.w1(32'h3b293163),
	.w2(32'h3bbbce93),
	.w3(32'h3beb731b),
	.w4(32'hbad435db),
	.w5(32'hbb21182a),
	.w6(32'hbaaf2be0),
	.w7(32'h3abbd76f),
	.w8(32'h3b32455f),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be20b17),
	.w1(32'hbcd5174b),
	.w2(32'hbd76880f),
	.w3(32'hbacced8c),
	.w4(32'hbc37c3a7),
	.w5(32'hbd230337),
	.w6(32'hbc2fe180),
	.w7(32'hbd060f36),
	.w8(32'hbca36b7c),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd55ffb2),
	.w1(32'hbc0aae91),
	.w2(32'hbd6c6be5),
	.w3(32'hbcf7148a),
	.w4(32'hbc54563b),
	.w5(32'hbd3cd4f9),
	.w6(32'hbb71acd8),
	.w7(32'hbca07621),
	.w8(32'hbcc617a9),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd63b818),
	.w1(32'h39d855bb),
	.w2(32'h3bb4645a),
	.w3(32'hbd0fe981),
	.w4(32'h3bac2da3),
	.w5(32'h3a9492c5),
	.w6(32'hba9cf5ca),
	.w7(32'h3bc0cd32),
	.w8(32'hb9c43bf5),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4106ec),
	.w1(32'hbbfe56e2),
	.w2(32'hbc724e39),
	.w3(32'hbb4e845c),
	.w4(32'hbbb945c3),
	.w5(32'h3acdeba3),
	.w6(32'hbbf8a42f),
	.w7(32'hbc467b82),
	.w8(32'hbc67e348),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc11abb6),
	.w1(32'hbc63663c),
	.w2(32'hbcca805c),
	.w3(32'hbb87b599),
	.w4(32'hbc15bcdd),
	.w5(32'hbcb76909),
	.w6(32'hbca1bd0e),
	.w7(32'hbcbca0af),
	.w8(32'hbc9c20a6),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc96694b),
	.w1(32'hbbdf1c67),
	.w2(32'hbba71fa3),
	.w3(32'hbc942efa),
	.w4(32'hbb43e5cd),
	.w5(32'hbb161ab8),
	.w6(32'hbbde6734),
	.w7(32'hbbdce120),
	.w8(32'hbc30ace8),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc197c57),
	.w1(32'hbb687025),
	.w2(32'hbab5bc3a),
	.w3(32'hbbdffa3e),
	.w4(32'hbb94a516),
	.w5(32'hba933f44),
	.w6(32'hbbd47a66),
	.w7(32'hbbe21762),
	.w8(32'hbbfef4bc),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf18f7e),
	.w1(32'hba916560),
	.w2(32'h3bc8015e),
	.w3(32'hbb55d55d),
	.w4(32'hbbb53844),
	.w5(32'h3aaf7cf9),
	.w6(32'hbb64838b),
	.w7(32'h3b4b6ae0),
	.w8(32'h3b52f0c6),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2b2cba),
	.w1(32'h3cc9128d),
	.w2(32'h3d2fdbcb),
	.w3(32'h3bb7695f),
	.w4(32'h3c7be25f),
	.w5(32'h3cb36578),
	.w6(32'h3c3af5e2),
	.w7(32'h3c7292fe),
	.w8(32'h3bed56b1),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca2c206),
	.w1(32'h3d0643f8),
	.w2(32'h3cd960fd),
	.w3(32'h3c721d2e),
	.w4(32'h3c80b3c6),
	.w5(32'h3c67505d),
	.w6(32'h3c8ed1eb),
	.w7(32'h3c48a4c5),
	.w8(32'h3b60f117),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb200fd),
	.w1(32'hbc12c519),
	.w2(32'hbd0c494d),
	.w3(32'h3c147995),
	.w4(32'hbc563f81),
	.w5(32'hbc9f1096),
	.w6(32'h392ade8c),
	.w7(32'hbcae12a0),
	.w8(32'hbc4dff61),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcdaa100),
	.w1(32'hbc823812),
	.w2(32'hbc9b1735),
	.w3(32'hbcd64b9c),
	.w4(32'hbb524a9f),
	.w5(32'hbc3086a5),
	.w6(32'hbbd9de9e),
	.w7(32'hbcbc7e1b),
	.w8(32'hbc65fc41),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc572630),
	.w1(32'hbc680d0b),
	.w2(32'hbbca07e6),
	.w3(32'hbc384b28),
	.w4(32'hbab5a531),
	.w5(32'hba45c46b),
	.w6(32'hbc180b52),
	.w7(32'hbc2cf562),
	.w8(32'hbc55e807),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb08e205),
	.w1(32'h3cf1a8cb),
	.w2(32'h3ca4f0c4),
	.w3(32'h3b74f756),
	.w4(32'h3c71e1bf),
	.w5(32'h3c85f9b1),
	.w6(32'h3c9ecde5),
	.w7(32'h3c8dcbb9),
	.w8(32'h3be372b1),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3befbb05),
	.w1(32'h3c1b877d),
	.w2(32'h3c844733),
	.w3(32'h3c49123e),
	.w4(32'hbb634db0),
	.w5(32'hbc0187f6),
	.w6(32'hbb95974e),
	.w7(32'h3b9b059d),
	.w8(32'h3bf19427),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadf793b),
	.w1(32'hbbeeedb8),
	.w2(32'hbb29a688),
	.w3(32'hbc2cd947),
	.w4(32'hbbbd7e4d),
	.w5(32'hbb0175d0),
	.w6(32'hbb321648),
	.w7(32'hba9e6e0c),
	.w8(32'hbadb23ad),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38815f71),
	.w1(32'hb9b5c80e),
	.w2(32'h3b59578e),
	.w3(32'hbb113458),
	.w4(32'h38bf5250),
	.w5(32'hbb201273),
	.w6(32'hbb9682ba),
	.w7(32'h3a844c02),
	.w8(32'h3b1762c0),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb4dc7c),
	.w1(32'hb9c48dcc),
	.w2(32'h3b3ae9c4),
	.w3(32'h3b0b1e27),
	.w4(32'h3ad65a6b),
	.w5(32'h3aef3598),
	.w6(32'h3c0cc9b3),
	.w7(32'h3c0fdf83),
	.w8(32'h3beb44d2),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae56c84),
	.w1(32'h3d025bef),
	.w2(32'h3cc34396),
	.w3(32'hbb149279),
	.w4(32'h3ccd9a4b),
	.w5(32'h3cdb8ba3),
	.w6(32'h3c5227c1),
	.w7(32'h3c9c6a5b),
	.w8(32'h3c0171c2),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf41ceb),
	.w1(32'hbce57ee5),
	.w2(32'hbda111a4),
	.w3(32'h3c2d594a),
	.w4(32'hbc74df13),
	.w5(32'hbd8441c7),
	.w6(32'hbbd047d1),
	.w7(32'hbcfa1e1a),
	.w8(32'hbccf127b),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd910410),
	.w1(32'hbcc333b6),
	.w2(32'hbd3f243b),
	.w3(32'hbd60086b),
	.w4(32'hbc4c9aa2),
	.w5(32'hbd1f0939),
	.w6(32'hbc4d6369),
	.w7(32'hbc92e923),
	.w8(32'hbc5eed5c),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd07f327),
	.w1(32'hb9fce4c7),
	.w2(32'h3ad0d717),
	.w3(32'hbd19e518),
	.w4(32'h3ae5a2aa),
	.w5(32'h3b840d27),
	.w6(32'hbb669170),
	.w7(32'hbb8f7784),
	.w8(32'hbb981772),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afcdc97),
	.w1(32'h3b83452d),
	.w2(32'h3bf3c921),
	.w3(32'h3a561c55),
	.w4(32'h3bb56ab7),
	.w5(32'h3c13ee69),
	.w6(32'h3b3f02e7),
	.w7(32'h3b8b4fe3),
	.w8(32'h3c1c9ba8),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c58abc5),
	.w1(32'hbcbf8611),
	.w2(32'hbce53c6b),
	.w3(32'h3c406e2f),
	.w4(32'hbc6070c4),
	.w5(32'hbc52271b),
	.w6(32'hbc0284c6),
	.w7(32'hbc9e662b),
	.w8(32'hbb5e4aa4),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc566f78),
	.w1(32'h3a6b48c7),
	.w2(32'hbaf6140c),
	.w3(32'hbc117e62),
	.w4(32'h3a1e5b81),
	.w5(32'hbaa637c3),
	.w6(32'hb90b2baf),
	.w7(32'hbb039846),
	.w8(32'hb9a995e1),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c905c7),
	.w1(32'hbac8847c),
	.w2(32'hbbe8a5d9),
	.w3(32'hbad851c7),
	.w4(32'h3c212cf0),
	.w5(32'h3bd62b15),
	.w6(32'hbbb57cc2),
	.w7(32'hbbdd9451),
	.w8(32'hbc2ec0a2),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b5a08),
	.w1(32'h3b010601),
	.w2(32'hbc58b813),
	.w3(32'hbc087294),
	.w4(32'h3b11c403),
	.w5(32'hbc3bece2),
	.w6(32'hbc59d4e0),
	.w7(32'hbc9f6a23),
	.w8(32'hbc880e28),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaa5e78),
	.w1(32'hbc17b260),
	.w2(32'hb903c340),
	.w3(32'hbc875ea8),
	.w4(32'hbb5a10ea),
	.w5(32'hbb417737),
	.w6(32'hbc491bee),
	.w7(32'hbc832e7f),
	.w8(32'hbc313676),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8113a5),
	.w1(32'hbb8e07e7),
	.w2(32'h3acf4e91),
	.w3(32'hbb168d09),
	.w4(32'hbbbb999f),
	.w5(32'h3a397751),
	.w6(32'hba96fcea),
	.w7(32'h3ade1458),
	.w8(32'hbc54d690),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf3c493),
	.w1(32'hbc308d68),
	.w2(32'h3b1c6b98),
	.w3(32'h3bfc4489),
	.w4(32'hbc047557),
	.w5(32'h3bac45ef),
	.w6(32'hbc5f083e),
	.w7(32'hbb708bcb),
	.w8(32'hbc01cfe3),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb02a688),
	.w1(32'h3ac4b840),
	.w2(32'h3a805e2b),
	.w3(32'hba3d8f9d),
	.w4(32'h3904cb9c),
	.w5(32'hbc1c9d66),
	.w6(32'h3afacc35),
	.w7(32'hbc0c9315),
	.w8(32'hbacb9181),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba5346d),
	.w1(32'hbce5d2a2),
	.w2(32'hbd89232a),
	.w3(32'hbbca8a20),
	.w4(32'hbca1f664),
	.w5(32'hbd633a44),
	.w6(32'hbcb872be),
	.w7(32'hbcf729b0),
	.w8(32'hbc947a33),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd5f80d3),
	.w1(32'h3b66d20e),
	.w2(32'hbb91d311),
	.w3(32'hbd5a91e1),
	.w4(32'h3c43e034),
	.w5(32'h3c08918b),
	.w6(32'h3b884876),
	.w7(32'hba23f286),
	.w8(32'h3a67b814),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b32b1d9),
	.w1(32'hbc7dc0cc),
	.w2(32'hbc923581),
	.w3(32'h3bc9bd5c),
	.w4(32'hbc5a7a0f),
	.w5(32'hbc93fe35),
	.w6(32'hbc9245d1),
	.w7(32'hbcb6d247),
	.w8(32'hbb378a36),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc653109),
	.w1(32'h3c138c54),
	.w2(32'hbab41c8e),
	.w3(32'hbbe05de4),
	.w4(32'h3a8ce0c6),
	.w5(32'hbbfb0545),
	.w6(32'h3b830ea7),
	.w7(32'hbb12eda1),
	.w8(32'hb99efb23),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5f4950),
	.w1(32'h3bd036db),
	.w2(32'h3c2bcf61),
	.w3(32'hbb8c8371),
	.w4(32'h3b7e5f60),
	.w5(32'h3c0f68e4),
	.w6(32'h3ba356eb),
	.w7(32'h3bdaad86),
	.w8(32'h3b196f9e),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a448c99),
	.w1(32'h3bc93797),
	.w2(32'hba848cea),
	.w3(32'hba9deb43),
	.w4(32'h38e9f3e3),
	.w5(32'h3c01aacd),
	.w6(32'hbb2a4135),
	.w7(32'hbb38a117),
	.w8(32'hbc6c07aa),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb566f79),
	.w1(32'hbcc45b33),
	.w2(32'hbd4a086f),
	.w3(32'h3ba97e84),
	.w4(32'hbcbe2263),
	.w5(32'hbd45562c),
	.w6(32'hbc52f014),
	.w7(32'hbcad5300),
	.w8(32'hbc508455),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd214ecb),
	.w1(32'hbc00b1f0),
	.w2(32'hbc4c9c2c),
	.w3(32'hbd0bbe1c),
	.w4(32'hbbe6b01a),
	.w5(32'hbc16b2a7),
	.w6(32'hbb9dcfe9),
	.w7(32'hbbe27345),
	.w8(32'hbbe90e76),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc292233),
	.w1(32'hbcdfb035),
	.w2(32'hbd6f7288),
	.w3(32'hbbdf6142),
	.w4(32'hbcbf374d),
	.w5(32'hbd7ec30e),
	.w6(32'hbc298853),
	.w7(32'hbcb6c715),
	.w8(32'hbc7a1ccf),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd435182),
	.w1(32'h3af8ab99),
	.w2(32'h3baca8bf),
	.w3(32'hbd4e8e80),
	.w4(32'hbb2249e9),
	.w5(32'hba9df7b6),
	.w6(32'h3ab9e4bf),
	.w7(32'hbb9d3bfc),
	.w8(32'hbabef103),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b36d353),
	.w1(32'h36c4cb2e),
	.w2(32'h3bdf62b0),
	.w3(32'h3accdcbf),
	.w4(32'hbb4a3170),
	.w5(32'hbb58df9a),
	.w6(32'hb9b7557e),
	.w7(32'h390e4457),
	.w8(32'h3ad48d96),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7b45d3),
	.w1(32'hb90232ff),
	.w2(32'hbc65afbe),
	.w3(32'h3b94d908),
	.w4(32'h3a8816d4),
	.w5(32'h3c1fe954),
	.w6(32'h3b8cbfe3),
	.w7(32'hbc4524ef),
	.w8(32'hbc87ad79),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc62c852),
	.w1(32'hb81f3498),
	.w2(32'h3b6fff30),
	.w3(32'h3b1b269a),
	.w4(32'h3b8e75e9),
	.w5(32'h3b06bb01),
	.w6(32'hba164a96),
	.w7(32'h397565ef),
	.w8(32'hbbb1401d),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac34574),
	.w1(32'hbaf2222c),
	.w2(32'h3a016d17),
	.w3(32'hbb97bc93),
	.w4(32'hb9a89caa),
	.w5(32'h3b7d6782),
	.w6(32'hba23d210),
	.w7(32'h39df36eb),
	.w8(32'hbac291b7),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb206b4b),
	.w1(32'h3c20ca62),
	.w2(32'h3c1e63f4),
	.w3(32'h3b100348),
	.w4(32'h3c92e2a8),
	.w5(32'h3ca3b7b8),
	.w6(32'h3b87d024),
	.w7(32'h3b2665f6),
	.w8(32'h3b613893),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4dcf01),
	.w1(32'h3b933bea),
	.w2(32'h3ba79a0f),
	.w3(32'h3ca85502),
	.w4(32'h3ac2faa4),
	.w5(32'h3c00ff4b),
	.w6(32'h3a893f86),
	.w7(32'h3b443f0e),
	.w8(32'h3a86a65b),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aac51fc),
	.w1(32'h3c9f8874),
	.w2(32'h3c93fbe3),
	.w3(32'h3b170185),
	.w4(32'h3bc29409),
	.w5(32'h3c645a8d),
	.w6(32'h3c721d1d),
	.w7(32'h3cb79fca),
	.w8(32'h3c0ece56),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7d2ebb),
	.w1(32'h3b3da2e6),
	.w2(32'hbae9f730),
	.w3(32'h3c0b5a80),
	.w4(32'h3aaa26b4),
	.w5(32'h39783ac5),
	.w6(32'hbb20a586),
	.w7(32'hb9f47575),
	.w8(32'hbbc10ddf),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc852e1),
	.w1(32'h3c788376),
	.w2(32'h3ce89131),
	.w3(32'hbbaa9881),
	.w4(32'h3c212fd4),
	.w5(32'h3c463158),
	.w6(32'h3c54f6c1),
	.w7(32'h3c9ffdeb),
	.w8(32'h3c1c8ebe),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc6f7b0),
	.w1(32'h3c131409),
	.w2(32'h3c76ed70),
	.w3(32'h3c2b5f76),
	.w4(32'h3c1497d3),
	.w5(32'h3c4229ae),
	.w6(32'h3b05716e),
	.w7(32'h3c81d7f6),
	.w8(32'h3c52531e),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4222cf),
	.w1(32'hbb2bb4d6),
	.w2(32'hbbd7c0e9),
	.w3(32'h3c2922b3),
	.w4(32'hbaa0153f),
	.w5(32'hbb037cc5),
	.w6(32'hbacdc518),
	.w7(32'hbb46a1a1),
	.w8(32'hba99ca96),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb38b169),
	.w1(32'h3b6cd491),
	.w2(32'h3bcbb7af),
	.w3(32'h3a228036),
	.w4(32'hbbd01bf9),
	.w5(32'h3b93523c),
	.w6(32'hbc03e639),
	.w7(32'hba8252ff),
	.w8(32'hbb9b4dbd),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baba05d),
	.w1(32'h3c3e4a46),
	.w2(32'h3bf5a099),
	.w3(32'h3ae49dee),
	.w4(32'h3c1177a8),
	.w5(32'h3c64415b),
	.w6(32'h3bfb6fa8),
	.w7(32'hbb8b46d6),
	.w8(32'h3ae0c923),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbda4216),
	.w1(32'h3b1d50e3),
	.w2(32'hbc8a9fcd),
	.w3(32'h3bb0c0b4),
	.w4(32'hbb959d78),
	.w5(32'hbc86ceff),
	.w6(32'hbab7f00d),
	.w7(32'h39bffa3e),
	.w8(32'hbb465c11),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9a03ff),
	.w1(32'hba367eca),
	.w2(32'h3ae59a67),
	.w3(32'hbc71cde6),
	.w4(32'h3a3913f2),
	.w5(32'h3a8c6b71),
	.w6(32'h3a47c97e),
	.w7(32'h3b12e32b),
	.w8(32'h3a3cb642),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad28e77),
	.w1(32'h3bcfc390),
	.w2(32'h3c675f46),
	.w3(32'hb9832697),
	.w4(32'hbb0b6beb),
	.w5(32'h3b701e29),
	.w6(32'h3c3cc8e8),
	.w7(32'h3c2477b6),
	.w8(32'hbb4c0175),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule