module layer_6_featuremap_72(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 2048;
	parameter IMG_SIZE = 52;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcce5ae8),
	.w1(32'h39b280d2),
	.w2(32'h3c045c83),
	.w3(32'hba5d3117),
	.w4(32'h3b4f4eea),
	.w5(32'hbbc5dd5c),
	.w6(32'h3b510a9e),
	.w7(32'h3c2b129a),
	.w8(32'h3a130705),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91472f0),
	.w1(32'hbbaa01e8),
	.w2(32'hbb5fc752),
	.w3(32'hba20109e),
	.w4(32'h3b32045f),
	.w5(32'h3bb73d9f),
	.w6(32'hbc14c5a6),
	.w7(32'hbbe44b76),
	.w8(32'h38ec4ba9),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b93eee1),
	.w1(32'hbb6c899f),
	.w2(32'hbc24bab6),
	.w3(32'hbb538b84),
	.w4(32'h3b6f3ce9),
	.w5(32'hbb329196),
	.w6(32'hbbd02ae5),
	.w7(32'hbc3d1a2b),
	.w8(32'hbb53d599),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbac6289),
	.w1(32'hbc5fbedd),
	.w2(32'hbc91f19c),
	.w3(32'hbc1f3590),
	.w4(32'hbc33870d),
	.w5(32'hbb04bcc9),
	.w6(32'hbc80527b),
	.w7(32'hbc9aa7c7),
	.w8(32'hbc107d01),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbec4eff),
	.w1(32'hbc5968dc),
	.w2(32'hbbf51c97),
	.w3(32'hbc126e02),
	.w4(32'hbbbbdc3a),
	.w5(32'h3836bee6),
	.w6(32'hbc0dac1e),
	.w7(32'hbb66387a),
	.w8(32'h3c21d31f),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c04d8f3),
	.w1(32'h3cfa487c),
	.w2(32'h3cf72f5c),
	.w3(32'h3cad3682),
	.w4(32'h3ca7e324),
	.w5(32'h3c4f47ca),
	.w6(32'h3d06ac6b),
	.w7(32'h3d09af75),
	.w8(32'h3cbe4a96),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca72103),
	.w1(32'hbd3241a9),
	.w2(32'hbd3275d1),
	.w3(32'hbd06e86b),
	.w4(32'hbd06e532),
	.w5(32'hbc452029),
	.w6(32'hbd4cc4f1),
	.w7(32'hbd51799f),
	.w8(32'hbcc73615),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc931782),
	.w1(32'hbc378fd5),
	.w2(32'hbc055dc2),
	.w3(32'hbc4bf827),
	.w4(32'hbbbf1827),
	.w5(32'hbc011045),
	.w6(32'hbc207a62),
	.w7(32'hbb3c9ddf),
	.w8(32'hbc59ca42),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7f96a1),
	.w1(32'h3bc42c56),
	.w2(32'hbb2cd109),
	.w3(32'hbbb904d5),
	.w4(32'h3ba9ccc8),
	.w5(32'h3c07f607),
	.w6(32'hbc28d532),
	.w7(32'h3af2f88a),
	.w8(32'h3b6bee6e),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc26f0dc),
	.w1(32'h3cd9b159),
	.w2(32'h3ccb4021),
	.w3(32'h3cbad130),
	.w4(32'h3cbae007),
	.w5(32'h3c0dc8d8),
	.w6(32'h3cf46e56),
	.w7(32'h3cf15f89),
	.w8(32'h3c5e7bc1),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c247c50),
	.w1(32'hbb37a0bf),
	.w2(32'hbbeb5d4b),
	.w3(32'h3909f66d),
	.w4(32'h3b323cea),
	.w5(32'hbc29d534),
	.w6(32'hbbdb4944),
	.w7(32'h3b894a93),
	.w8(32'hbabb14c6),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2b8ef4),
	.w1(32'hbb9fd264),
	.w2(32'hbb25853a),
	.w3(32'h39b3c64a),
	.w4(32'hbaee5f72),
	.w5(32'hbb92de43),
	.w6(32'hbb1c5f33),
	.w7(32'hbb0813f7),
	.w8(32'hba160865),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbec6a57),
	.w1(32'hbc185eec),
	.w2(32'hbbe3493c),
	.w3(32'hbb82b923),
	.w4(32'hbb4b00ab),
	.w5(32'hbb0dba61),
	.w6(32'hbbe9ae5e),
	.w7(32'hbb8db754),
	.w8(32'hbadee137),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc84119),
	.w1(32'hbb1514d1),
	.w2(32'hba4c8e21),
	.w3(32'hba50c901),
	.w4(32'hbb9e88f8),
	.w5(32'hbc3f9f62),
	.w6(32'hbb9bca3d),
	.w7(32'hbb4c2303),
	.w8(32'hbb78075f),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39eacefc),
	.w1(32'hbbec6009),
	.w2(32'hbb96ce2e),
	.w3(32'hba933a93),
	.w4(32'h3ba36128),
	.w5(32'h3c1259ac),
	.w6(32'hbbb885a1),
	.w7(32'hbb807787),
	.w8(32'h3a2f46e6),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a96033a),
	.w1(32'h3b70a626),
	.w2(32'h3c102c86),
	.w3(32'h3b4e3561),
	.w4(32'h3bb22c08),
	.w5(32'h3b105ae8),
	.w6(32'h3b2514af),
	.w7(32'h3bc48806),
	.w8(32'h3b734d0b),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b99c062),
	.w1(32'hbc2992ac),
	.w2(32'hbc41ecf4),
	.w3(32'hbc2bc69c),
	.w4(32'hbc190b5d),
	.w5(32'hbb9041b3),
	.w6(32'hbc01bdda),
	.w7(32'hbc0e222f),
	.w8(32'hba473068),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6b3231),
	.w1(32'h3bd9607e),
	.w2(32'h3c4bf436),
	.w3(32'h3bc50a09),
	.w4(32'h3c3a2cfa),
	.w5(32'h3a029e4e),
	.w6(32'h3c04d1b4),
	.w7(32'h3c5a3e36),
	.w8(32'h3a3b3382),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b10dd42),
	.w1(32'hbadbc0fe),
	.w2(32'hbbd0ea84),
	.w3(32'hbb9025e8),
	.w4(32'hbbca7084),
	.w5(32'hbb0ceca5),
	.w6(32'hbb4edf6b),
	.w7(32'hbbf4ecaf),
	.w8(32'hbbb582de),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb38b0c),
	.w1(32'h3b971d89),
	.w2(32'h3b952cc0),
	.w3(32'h3b389070),
	.w4(32'h379be69c),
	.w5(32'h3c03f594),
	.w6(32'h3ad7d1f9),
	.w7(32'h3bcf7bd9),
	.w8(32'h3c97893b),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c55ff3e),
	.w1(32'hbba0844a),
	.w2(32'hbbcedb12),
	.w3(32'hbb5ba164),
	.w4(32'hbb1cdf07),
	.w5(32'h3b425967),
	.w6(32'hbbee2985),
	.w7(32'hbc053346),
	.w8(32'hbb02d638),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8814c40),
	.w1(32'hbbbf2897),
	.w2(32'hbaf784e4),
	.w3(32'hba9c2826),
	.w4(32'h3a9cc71d),
	.w5(32'h3c135bf7),
	.w6(32'hbbdac78b),
	.w7(32'hbb337fc0),
	.w8(32'h3bba5a8b),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8c66f2),
	.w1(32'hbcaee675),
	.w2(32'hbcd03680),
	.w3(32'hbc29f749),
	.w4(32'hbc1d5634),
	.w5(32'hbc523e2e),
	.w6(32'hbc54d94e),
	.w7(32'hbc9769d1),
	.w8(32'hbcd8217e),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcfdd2a6),
	.w1(32'h3c5fc464),
	.w2(32'h3c460d9c),
	.w3(32'h3bb03e31),
	.w4(32'h3b61967d),
	.w5(32'h3b52371b),
	.w6(32'h3be686ea),
	.w7(32'h3b995770),
	.w8(32'h38e2d85f),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af4636f),
	.w1(32'hbb3b8f3c),
	.w2(32'hba42f9c6),
	.w3(32'hbbce2c19),
	.w4(32'h3a22a436),
	.w5(32'h3bc5eac6),
	.w6(32'hbbec00a9),
	.w7(32'h3b32b377),
	.w8(32'h3c364c71),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb092b07),
	.w1(32'h3b0c42f2),
	.w2(32'h3c038729),
	.w3(32'h3b68ca37),
	.w4(32'h3b816f21),
	.w5(32'h3bee48cc),
	.w6(32'h3b655616),
	.w7(32'h3c2a777f),
	.w8(32'h3bf73fc7),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c066a0b),
	.w1(32'hbb3fe23e),
	.w2(32'hbaec9830),
	.w3(32'hbadd8983),
	.w4(32'hbb7057c8),
	.w5(32'hbb1ef51b),
	.w6(32'hbbb0b585),
	.w7(32'hbb567e15),
	.w8(32'hba84f031),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba96323a),
	.w1(32'hbcc225a7),
	.w2(32'hbcce16cf),
	.w3(32'hbcb47224),
	.w4(32'hbca49ae1),
	.w5(32'hb97479f5),
	.w6(32'hbcf1f1d9),
	.w7(32'hbcfd8360),
	.w8(32'hbc1984f4),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba19c54),
	.w1(32'hbb7cd0ec),
	.w2(32'hbb9bc3d2),
	.w3(32'hb9962a7b),
	.w4(32'hba522ac1),
	.w5(32'hbaf5ab4f),
	.w6(32'hbb3e82b3),
	.w7(32'hbb5d5cc3),
	.w8(32'hbb87f17e),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc097693),
	.w1(32'h3b92c279),
	.w2(32'h3c1c28a1),
	.w3(32'hbb873699),
	.w4(32'h3c1c65db),
	.w5(32'h3c3c1e85),
	.w6(32'hbb27005a),
	.w7(32'h3c15d29a),
	.w8(32'h3c7b68e5),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4d6a6a),
	.w1(32'hbbd8f5e1),
	.w2(32'hbacbf116),
	.w3(32'hbb55a69d),
	.w4(32'hbbcdda74),
	.w5(32'hbc10b27a),
	.w6(32'hbbde8097),
	.w7(32'hbc34fe6e),
	.w8(32'hbc365477),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba4941a),
	.w1(32'hba567bb5),
	.w2(32'h3c33cf71),
	.w3(32'h3ad5041c),
	.w4(32'h3bb16d75),
	.w5(32'hbbb04db8),
	.w6(32'h3c36be39),
	.w7(32'h3c9fea47),
	.w8(32'h3bacbfaa),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1fbddf),
	.w1(32'h3bbf9d24),
	.w2(32'h3a84b414),
	.w3(32'h3b4e04ba),
	.w4(32'h3c4402a5),
	.w5(32'h3c61c6ed),
	.w6(32'h3baef614),
	.w7(32'h3b9df290),
	.w8(32'h3cc4e671),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c86f087),
	.w1(32'h3b639dfb),
	.w2(32'h3bdd7ac4),
	.w3(32'hbb86618f),
	.w4(32'h3ac9700b),
	.w5(32'h3b68dfe0),
	.w6(32'h3b28ee0a),
	.w7(32'h39e33637),
	.w8(32'h3c684ac9),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5045aa),
	.w1(32'h3c5c0624),
	.w2(32'h3bc6bedf),
	.w3(32'h3c129f96),
	.w4(32'h3b436f73),
	.w5(32'hbb498b6d),
	.w6(32'h3c5fe32f),
	.w7(32'h3bd73579),
	.w8(32'h3a00ff53),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2a591c),
	.w1(32'hbbb5afb2),
	.w2(32'h3a1bb1c9),
	.w3(32'hb9d9d765),
	.w4(32'hbb27386b),
	.w5(32'h3b0f52cf),
	.w6(32'h3b3c2c12),
	.w7(32'hba038691),
	.w8(32'h3c238b8c),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba34aba),
	.w1(32'h3b40f8f1),
	.w2(32'h3c3a8a0c),
	.w3(32'hba97f9a2),
	.w4(32'h3b484d53),
	.w5(32'hbb86ff01),
	.w6(32'h3be704e2),
	.w7(32'h3c6b0b79),
	.w8(32'h3ba6a47a),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9c7d8a),
	.w1(32'hbc4d3062),
	.w2(32'hbbe7ce9e),
	.w3(32'hbc136622),
	.w4(32'hbba81d87),
	.w5(32'hb773f3c9),
	.w6(32'hbc4ae066),
	.w7(32'hbc09a6f1),
	.w8(32'hbb496748),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2c8366),
	.w1(32'hba5b539e),
	.w2(32'hbae01614),
	.w3(32'hba2ddff6),
	.w4(32'h3adcdc22),
	.w5(32'hbbf5a59c),
	.w6(32'hbb9f51b5),
	.w7(32'hbc216358),
	.w8(32'hbc30b004),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc79c63d),
	.w1(32'hba2aac66),
	.w2(32'hbb869c59),
	.w3(32'hbb1111ae),
	.w4(32'hba32ce6e),
	.w5(32'hba85169b),
	.w6(32'hbc56c6b4),
	.w7(32'h39fc03a1),
	.w8(32'h3a9502ec),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8acbae),
	.w1(32'h3bd59a05),
	.w2(32'hba8e4eb0),
	.w3(32'hbb8d2b7f),
	.w4(32'h3ae1763e),
	.w5(32'hbbb50bc4),
	.w6(32'h3a59bb16),
	.w7(32'h3bc1d1c7),
	.w8(32'h3a5550cc),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b32b881),
	.w1(32'hbc591cfe),
	.w2(32'hbc8b38a1),
	.w3(32'hbc30f478),
	.w4(32'hbc45bd3a),
	.w5(32'hbb0ea7c6),
	.w6(32'hbc83bd7b),
	.w7(32'hbc9fb16f),
	.w8(32'hbbe6431c),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcd5186),
	.w1(32'h3b8d46ca),
	.w2(32'h3c1efee9),
	.w3(32'h3ba7f687),
	.w4(32'h3c1da92f),
	.w5(32'h3bf17d47),
	.w6(32'h3bf65bf5),
	.w7(32'h3c6c1f7a),
	.w8(32'h3bf8488e),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b696005),
	.w1(32'hbbdb6617),
	.w2(32'hbb411aa8),
	.w3(32'h3ad570df),
	.w4(32'hbac2f7a1),
	.w5(32'h3c5bfc0a),
	.w6(32'hba0b7fbc),
	.w7(32'hb9b59822),
	.w8(32'h3c395b1b),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b13ab1c),
	.w1(32'hbbf686e6),
	.w2(32'hbbdf19c8),
	.w3(32'hbbb15018),
	.w4(32'hbb65fc8e),
	.w5(32'hba8423f2),
	.w6(32'hbbdcc000),
	.w7(32'hbbb0e4b0),
	.w8(32'hbb179d94),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6210c9),
	.w1(32'hbc55f0f5),
	.w2(32'hbc15fec3),
	.w3(32'h3c29fddd),
	.w4(32'h3c476e92),
	.w5(32'h3b79700b),
	.w6(32'hb8bfb301),
	.w7(32'h3aec7a32),
	.w8(32'h3b8ef0b2),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb225b0c),
	.w1(32'hbbcb5609),
	.w2(32'hbc590128),
	.w3(32'h3b020f8b),
	.w4(32'hba290043),
	.w5(32'h3c90a1d3),
	.w6(32'h3a8d3ea8),
	.w7(32'hbc1336ca),
	.w8(32'h3c51f9c3),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c623c51),
	.w1(32'h3ad2076c),
	.w2(32'h3ca3ed2b),
	.w3(32'hbbbcd506),
	.w4(32'h3c31a99f),
	.w5(32'h3c38b8d5),
	.w6(32'hbbcadfc0),
	.w7(32'h3c8b16d3),
	.w8(32'h3c9d22df),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8a32d0),
	.w1(32'h3afc5a24),
	.w2(32'hb90ff0bf),
	.w3(32'h3b3e6c8c),
	.w4(32'h3b21e296),
	.w5(32'h3bb2e0cd),
	.w6(32'h3a95e2ec),
	.w7(32'h37e16294),
	.w8(32'h3b70ed2c),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4d0537),
	.w1(32'hbc32039d),
	.w2(32'h3bc82f4d),
	.w3(32'h3c122dd8),
	.w4(32'hbb9e4388),
	.w5(32'hbc593810),
	.w6(32'h3b0f0d3e),
	.w7(32'hbbb0512d),
	.w8(32'h3ba9d768),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8b843f),
	.w1(32'hbc34660f),
	.w2(32'hbcd2d604),
	.w3(32'hbb33631f),
	.w4(32'hbc6879cf),
	.w5(32'h3b90a447),
	.w6(32'hbc41d2dd),
	.w7(32'hbce0fcab),
	.w8(32'hbbb25bbf),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb37763),
	.w1(32'hbbd563a6),
	.w2(32'hbc797795),
	.w3(32'hbb8b53a5),
	.w4(32'hbc3bc90b),
	.w5(32'h3a2cd74f),
	.w6(32'hbc2b323f),
	.w7(32'hbca54503),
	.w8(32'hbbc9be23),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb619e6b),
	.w1(32'hbc70e55f),
	.w2(32'hbcaec7f7),
	.w3(32'hbc04dc65),
	.w4(32'hbc0f071d),
	.w5(32'h3beed01e),
	.w6(32'hbc9752da),
	.w7(32'hbcc4be12),
	.w8(32'hbbee0aa2),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd081a2),
	.w1(32'hbd31b2f0),
	.w2(32'hbd3404d4),
	.w3(32'hbcf366b1),
	.w4(32'hbccff0e0),
	.w5(32'hbba488f1),
	.w6(32'hbd3d8e51),
	.w7(32'hbd3c7021),
	.w8(32'hbcc13059),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc16dd1),
	.w1(32'hbc5daa72),
	.w2(32'hbcbee97c),
	.w3(32'hbb014d68),
	.w4(32'hbc09fc12),
	.w5(32'h3b009842),
	.w6(32'hbc823560),
	.w7(32'hbcbf167e),
	.w8(32'hbc111dc6),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc42fbe0),
	.w1(32'h3b23bfa3),
	.w2(32'hbaef3df8),
	.w3(32'hbbec3f48),
	.w4(32'hbba6fbc0),
	.w5(32'hbaa4eb5b),
	.w6(32'hbb6d5924),
	.w7(32'hbc4cbd46),
	.w8(32'hbc3d47ba),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b05d549),
	.w1(32'h3b5cc03a),
	.w2(32'h3c04861e),
	.w3(32'h3bcf76d6),
	.w4(32'h3c00507c),
	.w5(32'h3c2c4ac4),
	.w6(32'h3c0916be),
	.w7(32'h3c5ec7b9),
	.w8(32'h3ca5e3c6),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0f4579),
	.w1(32'h3b3f4265),
	.w2(32'h3c029188),
	.w3(32'h3b4531ae),
	.w4(32'hbb3c4123),
	.w5(32'hba4dae7b),
	.w6(32'h3c0e105a),
	.w7(32'hba271354),
	.w8(32'hbbde8177),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf2f43e),
	.w1(32'hb99cc950),
	.w2(32'hbb3e2afe),
	.w3(32'hbb6f3ede),
	.w4(32'hbb98d33b),
	.w5(32'hbbc6d368),
	.w6(32'hbae912df),
	.w7(32'hbb99266e),
	.w8(32'hbbd93615),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1ed74f),
	.w1(32'hbabd1020),
	.w2(32'h3bcc5090),
	.w3(32'h3a10c811),
	.w4(32'hbb0db537),
	.w5(32'h3bbe0745),
	.w6(32'h3c23f539),
	.w7(32'h3bbb9c82),
	.w8(32'h3cad6c7e),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4bacb8),
	.w1(32'hbbe6a882),
	.w2(32'hbc2a64ca),
	.w3(32'hbc1741fc),
	.w4(32'hbc4e02d9),
	.w5(32'hbc67558e),
	.w6(32'hbc23b774),
	.w7(32'hbc5573f6),
	.w8(32'hbc973db5),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc38a01e),
	.w1(32'h3ab6a296),
	.w2(32'h3a156440),
	.w3(32'hbb1cfc6f),
	.w4(32'hbb9ac194),
	.w5(32'hbae867e8),
	.w6(32'h3b2dd4dd),
	.w7(32'hb9704e0c),
	.w8(32'hbb81af6b),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395b7110),
	.w1(32'h3b974ddd),
	.w2(32'hb9c1566e),
	.w3(32'hbc0f1f31),
	.w4(32'h3a7a532b),
	.w5(32'h3ba36326),
	.w6(32'hbc592dd9),
	.w7(32'hbc0686c1),
	.w8(32'h3c95a255),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bee49c9),
	.w1(32'h3c1f4acb),
	.w2(32'hbaa358c9),
	.w3(32'hbba36ca6),
	.w4(32'hbc984cc9),
	.w5(32'hbce6582d),
	.w6(32'h3b91b70d),
	.w7(32'hbc3e5f82),
	.w8(32'hbcd663c6),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

endmodule