module layer_8_featuremap_214(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2a615f),
	.w1(32'h3bc5c91c),
	.w2(32'h3cfc3ac8),
	.w3(32'h3bfb99e0),
	.w4(32'h383a717a),
	.w5(32'h3c8fc8c2),
	.w6(32'h3c3013a9),
	.w7(32'h3cc79481),
	.w8(32'h3c9f2874),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc70e83),
	.w1(32'h381e7f3d),
	.w2(32'hba4a7810),
	.w3(32'h3c6c394a),
	.w4(32'hbbf87f3a),
	.w5(32'hbc10e654),
	.w6(32'hb8164d10),
	.w7(32'h3ba0b2a4),
	.w8(32'h3b3c37fa),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9c4dda),
	.w1(32'h3c17021b),
	.w2(32'h3bc04f6a),
	.w3(32'h3acde540),
	.w4(32'hbba7a907),
	.w5(32'hbc47b7ce),
	.w6(32'h3b5bf158),
	.w7(32'h3ba6480c),
	.w8(32'h3b82b676),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e1a26),
	.w1(32'hbc777ec5),
	.w2(32'hbbc38a3c),
	.w3(32'hbbbd065c),
	.w4(32'hbc079903),
	.w5(32'hbb76d7a4),
	.w6(32'h3c06d906),
	.w7(32'h3c218f06),
	.w8(32'h3c14e63c),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b77b5),
	.w1(32'h3afad75c),
	.w2(32'h3a89405c),
	.w3(32'hbc2f03f4),
	.w4(32'h3bf79825),
	.w5(32'h3c0080a8),
	.w6(32'hbb175675),
	.w7(32'hbbfb8035),
	.w8(32'hbbfabf79),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b963eed),
	.w1(32'hbae93693),
	.w2(32'hbc72167c),
	.w3(32'h3c375458),
	.w4(32'hbc92cbe7),
	.w5(32'hbd172d25),
	.w6(32'hbb70819f),
	.w7(32'hbc798980),
	.w8(32'hbc8284e6),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb479b9e),
	.w1(32'h3a454348),
	.w2(32'hbb361328),
	.w3(32'hbc1f875a),
	.w4(32'h3c1b5c1f),
	.w5(32'h3c1f2659),
	.w6(32'hbbad3e2f),
	.w7(32'hbc27a56a),
	.w8(32'hbc370fcd),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc81aa10),
	.w1(32'hbbe5b843),
	.w2(32'h3bf18356),
	.w3(32'hba3c2d75),
	.w4(32'hbc2c7e17),
	.w5(32'hbc073941),
	.w6(32'hba024cfc),
	.w7(32'h3c1c763f),
	.w8(32'h3c289cc4),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be7bc24),
	.w1(32'hbb8acf2a),
	.w2(32'hbb50c0f9),
	.w3(32'hbb5fed5f),
	.w4(32'hbc494005),
	.w5(32'hbc5812e1),
	.w6(32'h3a3465fe),
	.w7(32'h3af6edf7),
	.w8(32'hb9e3ba70),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb61599),
	.w1(32'h3a1d051c),
	.w2(32'h3ca3e174),
	.w3(32'hbc8b1ce6),
	.w4(32'h3c05b26c),
	.w5(32'h3c6e4639),
	.w6(32'h3b1ea8c6),
	.w7(32'h3c5a2f1e),
	.w8(32'h3c2a6daa),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfe3d44),
	.w1(32'hbc5ee136),
	.w2(32'hbbc19a30),
	.w3(32'h3c237d57),
	.w4(32'hbc304428),
	.w5(32'hbb350f8f),
	.w6(32'hb91afc00),
	.w7(32'h3c017476),
	.w8(32'h3c2aa60d),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce7002a),
	.w1(32'hbc82be03),
	.w2(32'hbb97a90d),
	.w3(32'hbc635a88),
	.w4(32'h3bbbcb11),
	.w5(32'h3c2ab845),
	.w6(32'h3790386c),
	.w7(32'h3be295a5),
	.w8(32'hbb088a38),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4e99d0),
	.w1(32'h3ae6b73e),
	.w2(32'h3bb8f925),
	.w3(32'h3b39302b),
	.w4(32'h3b251032),
	.w5(32'hbc6fed31),
	.w6(32'h3afdc5da),
	.w7(32'h3b991134),
	.w8(32'h3a8d59de),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb1bfdd),
	.w1(32'h3b758e36),
	.w2(32'h3af84220),
	.w3(32'hbb0b54d7),
	.w4(32'h3a15f69f),
	.w5(32'hbbaea420),
	.w6(32'h3b95707e),
	.w7(32'hbb812c6c),
	.w8(32'hb995b5b7),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba7c0ad),
	.w1(32'hbae8d6c3),
	.w2(32'hbb33b37b),
	.w3(32'hb847491b),
	.w4(32'h3983aa62),
	.w5(32'hba4337f4),
	.w6(32'hbac6f319),
	.w7(32'hbb82e0e9),
	.w8(32'hbaa87b42),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa444fa),
	.w1(32'hbbb51040),
	.w2(32'h3b02f75c),
	.w3(32'hba12a872),
	.w4(32'hbca07b6b),
	.w5(32'hbb92b3ab),
	.w6(32'h3b9e4774),
	.w7(32'h3c59d598),
	.w8(32'h3c16938b),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3087f7),
	.w1(32'hbb976d6c),
	.w2(32'hbb2acea4),
	.w3(32'h3b9d86bb),
	.w4(32'hbc81b355),
	.w5(32'hb99af0d4),
	.w6(32'hba76c623),
	.w7(32'hbb5d63c6),
	.w8(32'h3bd47d51),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8aee8d),
	.w1(32'hbbaa741c),
	.w2(32'h3b22f989),
	.w3(32'h3bbd0e44),
	.w4(32'hbbe752c1),
	.w5(32'hbbb69aa7),
	.w6(32'h3bde7f2e),
	.w7(32'h3cc86cd4),
	.w8(32'h3c23c95c),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd54b980),
	.w1(32'hbd0b3196),
	.w2(32'h3c204bf0),
	.w3(32'h3c4833e7),
	.w4(32'h3b741a2b),
	.w5(32'h3d2047cd),
	.w6(32'h3c4e8e1e),
	.w7(32'h3d53acb3),
	.w8(32'h3cf564c1),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c85a1b4),
	.w1(32'h3b8a6a66),
	.w2(32'hbaa75685),
	.w3(32'h3abe8e41),
	.w4(32'h3b3ac9bc),
	.w5(32'hbbae3509),
	.w6(32'hbbdbdebe),
	.w7(32'hbb21b574),
	.w8(32'hbbfe5b8d),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfdeba2),
	.w1(32'hba9b8628),
	.w2(32'hbc7a7b9c),
	.w3(32'h3c1ef42f),
	.w4(32'hbc599246),
	.w5(32'hbcaecf29),
	.w6(32'hbbc18f6c),
	.w7(32'hbba14439),
	.w8(32'hbb7d1465),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe17895),
	.w1(32'h3b86db8a),
	.w2(32'h3c3559a2),
	.w3(32'hbc199836),
	.w4(32'hbad61d95),
	.w5(32'h3b298106),
	.w6(32'hbc05c6ab),
	.w7(32'hbb84e4aa),
	.w8(32'hbc4dab36),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd134be5),
	.w1(32'hbd2195e0),
	.w2(32'h3c8e9f50),
	.w3(32'hbc5d5bbb),
	.w4(32'hbcf59fba),
	.w5(32'h3b9a88d1),
	.w6(32'h3b2c1536),
	.w7(32'h3cdfcf91),
	.w8(32'h3d250c36),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c159d7c),
	.w1(32'h3c1152fd),
	.w2(32'h3ae7fb1e),
	.w3(32'hbbada1e4),
	.w4(32'h3a21ee43),
	.w5(32'h3a485b86),
	.w6(32'hbbced53c),
	.w7(32'hbad2c858),
	.w8(32'hbbe8c5d5),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb006d6c),
	.w1(32'h3b1422b7),
	.w2(32'h3b498274),
	.w3(32'h3b01fc9f),
	.w4(32'hbb3b0ee5),
	.w5(32'hba70b57c),
	.w6(32'h3bccf810),
	.w7(32'hba0a7915),
	.w8(32'h3aabc3b6),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc26fe34),
	.w1(32'h3b2d1ea8),
	.w2(32'h3cf174a6),
	.w3(32'h3af1d92b),
	.w4(32'h3c2e7687),
	.w5(32'h3c5e4572),
	.w6(32'h3c95ece5),
	.w7(32'h3cbfcfa6),
	.w8(32'h3c76de70),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cf720e2),
	.w1(32'hbbc9eb49),
	.w2(32'hbba69471),
	.w3(32'h3c8d5bc6),
	.w4(32'hbc97264c),
	.w5(32'hbc31c265),
	.w6(32'hbb286607),
	.w7(32'h3a2a5f90),
	.w8(32'h3b80128b),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd9ad442),
	.w1(32'hbd6b6517),
	.w2(32'hbd1123e3),
	.w3(32'h3c9bb646),
	.w4(32'hbd740da1),
	.w5(32'hbd553887),
	.w6(32'h3cc4ce3c),
	.w7(32'h3d46367a),
	.w8(32'h3cc998db),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc96635b),
	.w1(32'hbb2e7cfc),
	.w2(32'h3c14cba7),
	.w3(32'hbc384a7b),
	.w4(32'h3bcd40c1),
	.w5(32'h3bef322a),
	.w6(32'h3a0a50f8),
	.w7(32'h3c8c69ec),
	.w8(32'h3c5cc4d6),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac3b710),
	.w1(32'hb9b78422),
	.w2(32'hbb895fd3),
	.w3(32'hbbbec725),
	.w4(32'h3bb98ec1),
	.w5(32'h3c077bee),
	.w6(32'hbb8f19a5),
	.w7(32'hbbb26614),
	.w8(32'hbb6350a9),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1c68c7),
	.w1(32'hbb34d83e),
	.w2(32'h3ac848b0),
	.w3(32'h3c419dde),
	.w4(32'h3aa01806),
	.w5(32'h3b9c13a7),
	.w6(32'hbb9a8490),
	.w7(32'hbb20878f),
	.w8(32'h3b5773fd),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf0f3e1),
	.w1(32'h3bf7e3b8),
	.w2(32'h3b539eb8),
	.w3(32'h3a72c47b),
	.w4(32'hb90d4b8d),
	.w5(32'h3b347405),
	.w6(32'hb9b02fa7),
	.w7(32'hbad74fb1),
	.w8(32'h3abbb480),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b861874),
	.w1(32'h3acf9168),
	.w2(32'hbaa966bc),
	.w3(32'h3c08d0cc),
	.w4(32'hbca41034),
	.w5(32'hbc604a46),
	.w6(32'h3c17ea3d),
	.w7(32'h3caf2036),
	.w8(32'h3c2634b3),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3befc78c),
	.w1(32'hbb8144c1),
	.w2(32'hbb2b95c0),
	.w3(32'hbc164cd6),
	.w4(32'h3b270776),
	.w5(32'h3c60e473),
	.w6(32'hbba23766),
	.w7(32'hbbe4ebaa),
	.w8(32'hbbcbefb3),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad1da70),
	.w1(32'hbb997bca),
	.w2(32'hbba663c7),
	.w3(32'h3b8bb76d),
	.w4(32'hbc6a374e),
	.w5(32'hbc8d9b49),
	.w6(32'hbc764536),
	.w7(32'hbc273f5a),
	.w8(32'hbbb44a2c),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3d7d74),
	.w1(32'hbccea8b8),
	.w2(32'hbcbd1b1d),
	.w3(32'hbc0291f2),
	.w4(32'h3a1f934c),
	.w5(32'h3b8344c1),
	.w6(32'hbc355680),
	.w7(32'hbbcb195c),
	.w8(32'hbc00c948),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5ed21b),
	.w1(32'h3924124c),
	.w2(32'h3a93b293),
	.w3(32'h3b88cd43),
	.w4(32'hbb511064),
	.w5(32'h377e09e0),
	.w6(32'h3a7d6667),
	.w7(32'h3b5d3bb5),
	.w8(32'h3b47a48e),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa8515b),
	.w1(32'hbba5f84c),
	.w2(32'hbbc94e15),
	.w3(32'hbb2d452b),
	.w4(32'hbbea9771),
	.w5(32'hbc1a07ed),
	.w6(32'h3ada1705),
	.w7(32'h3ab7b443),
	.w8(32'h3be19f2a),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9c0f90),
	.w1(32'h3ac7ab1a),
	.w2(32'h3b7ce0fa),
	.w3(32'hbb39be20),
	.w4(32'hb9acc395),
	.w5(32'h3bcf484d),
	.w6(32'hbbba0021),
	.w7(32'hbb82d0d9),
	.w8(32'hbc0a6b30),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb382b46),
	.w1(32'hbb2538a7),
	.w2(32'hbba89842),
	.w3(32'h3be780a9),
	.w4(32'h3bf05405),
	.w5(32'h3c8ec623),
	.w6(32'hbb8622a1),
	.w7(32'hbc522caa),
	.w8(32'hbc0ad124),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd306bc0),
	.w1(32'hbc561f37),
	.w2(32'h3bdacb89),
	.w3(32'hbc54a146),
	.w4(32'h3c03830b),
	.w5(32'h3b0d0af5),
	.w6(32'h3c7404e4),
	.w7(32'h3d3adb94),
	.w8(32'h3cd511a2),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2bb9ad),
	.w1(32'hbbfde7e8),
	.w2(32'hbb7b17ad),
	.w3(32'hbb877a9d),
	.w4(32'hbc9a555c),
	.w5(32'hba9b5fc6),
	.w6(32'h39f71e8d),
	.w7(32'hbb1e293f),
	.w8(32'hbac29630),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8790aeb),
	.w1(32'h3bb768a6),
	.w2(32'h3b05b070),
	.w3(32'h3a9da537),
	.w4(32'h3a209d78),
	.w5(32'h3b20a1da),
	.w6(32'h3b9e7ab8),
	.w7(32'h3b9ad7d3),
	.w8(32'h3b8bf03d),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb844ce9),
	.w1(32'hbc1c7cdd),
	.w2(32'h3a0222e3),
	.w3(32'hbb075c63),
	.w4(32'hbbe4404c),
	.w5(32'h3b66ba74),
	.w6(32'hbb2c19bf),
	.w7(32'h3bbe83b4),
	.w8(32'h3ba78015),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc99b612),
	.w1(32'hbca8dcdb),
	.w2(32'h3baa48bb),
	.w3(32'h3b7b1904),
	.w4(32'hbc7cc52b),
	.w5(32'hbb18fc3a),
	.w6(32'h3bbd976f),
	.w7(32'h3cc96562),
	.w8(32'h3d08f5bf),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb96b73b),
	.w1(32'hbc26c128),
	.w2(32'h3a943ab1),
	.w3(32'hbbb5ec18),
	.w4(32'hba978a0e),
	.w5(32'h3c121e2d),
	.w6(32'hbabf64c6),
	.w7(32'hb99fc1c4),
	.w8(32'h39e2def1),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba6216d),
	.w1(32'h3b9ec45a),
	.w2(32'h3ba85b55),
	.w3(32'h3b2d9076),
	.w4(32'h3ce03f4b),
	.w5(32'h3d120e8f),
	.w6(32'hbc84c4a8),
	.w7(32'hbcc2e684),
	.w8(32'hbccc8b59),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc903934),
	.w1(32'hbc9740c9),
	.w2(32'h3b912e62),
	.w3(32'h3cb4b0ef),
	.w4(32'hbc1be31b),
	.w5(32'h3aea1236),
	.w6(32'hbbb04afd),
	.w7(32'h3b3ceb90),
	.w8(32'h3c70fe65),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2b1542),
	.w1(32'h3b6d750f),
	.w2(32'h3b9c2ee2),
	.w3(32'h3a4fe4e9),
	.w4(32'hbbe5dac3),
	.w5(32'hbbaea315),
	.w6(32'h3b1e995f),
	.w7(32'h3bbe8976),
	.w8(32'h3abfa2eb),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1ecb20),
	.w1(32'hbba49bc5),
	.w2(32'h3c00d01e),
	.w3(32'hbc3cc7c5),
	.w4(32'hbc19eb60),
	.w5(32'h3b55c158),
	.w6(32'h3c26ff6d),
	.w7(32'h3d060ef5),
	.w8(32'h3ccf16db),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be555f8),
	.w1(32'hbb0bb81a),
	.w2(32'hba7abd33),
	.w3(32'hbc14c806),
	.w4(32'hb9ec8b39),
	.w5(32'h3b6f036b),
	.w6(32'hbbf0ef8a),
	.w7(32'hba96d2e7),
	.w8(32'hbc28edd2),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd4b066),
	.w1(32'hbc5357b0),
	.w2(32'h3b87a230),
	.w3(32'hbc2f9946),
	.w4(32'hbcac8ad6),
	.w5(32'h3b9e513e),
	.w6(32'h3cb24251),
	.w7(32'h3d1445f2),
	.w8(32'h3d076cec),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafb5842),
	.w1(32'hbb69f4f2),
	.w2(32'h39ef38e3),
	.w3(32'hbbb5969a),
	.w4(32'hba9b366b),
	.w5(32'h3b9ee08d),
	.w6(32'h3aa7447d),
	.w7(32'h3bf4d54a),
	.w8(32'h3bcb2eb3),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3e1476),
	.w1(32'hbcbb78c7),
	.w2(32'hbbdf90fb),
	.w3(32'hbb948f55),
	.w4(32'h3b2e2aa3),
	.w5(32'h3b46b9d2),
	.w6(32'hbc76b0d9),
	.w7(32'h3c2bb029),
	.w8(32'h3c578e90),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb94820f),
	.w1(32'h3b0eb842),
	.w2(32'h3c0c4358),
	.w3(32'hbb94c851),
	.w4(32'hbc3205e6),
	.w5(32'hbc28993e),
	.w6(32'h3c205438),
	.w7(32'h3c8edbc3),
	.w8(32'h3c5d94f8),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5ef6c6),
	.w1(32'hbd1ec9e2),
	.w2(32'hbaf1454a),
	.w3(32'hbbac6a91),
	.w4(32'hbb32eb0f),
	.w5(32'h3c82417d),
	.w6(32'hbcb1b235),
	.w7(32'hbbec78ca),
	.w8(32'hbb08c44d),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2a8444),
	.w1(32'hbc0c1dc7),
	.w2(32'hba2e780b),
	.w3(32'h3b2b252d),
	.w4(32'hbc9f978b),
	.w5(32'hbcacb9f5),
	.w6(32'hbbe3b5e5),
	.w7(32'h3ae9baea),
	.w8(32'h3ba32fec),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb305573),
	.w1(32'hbc093270),
	.w2(32'hbb4e39a7),
	.w3(32'hbc67a1aa),
	.w4(32'hbc2d8eb5),
	.w5(32'hbb9d5259),
	.w6(32'h3b5429ff),
	.w7(32'h3b9a714b),
	.w8(32'h3b6dd7eb),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe643c6),
	.w1(32'hbc074244),
	.w2(32'hbb0b9125),
	.w3(32'hbc27c915),
	.w4(32'hbbb70a9e),
	.w5(32'h3a9d2acd),
	.w6(32'hba84e57c),
	.w7(32'h3aaf49b6),
	.w8(32'h3c0335a0),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb56953),
	.w1(32'hba4fdb8c),
	.w2(32'h3b39ab65),
	.w3(32'h3958e93f),
	.w4(32'h3b0c6c2e),
	.w5(32'h3beeb99f),
	.w6(32'h3b7c4a95),
	.w7(32'h3c631c3e),
	.w8(32'h3c3a9811),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b31c427),
	.w1(32'hba88f358),
	.w2(32'h3b479875),
	.w3(32'h3a4f5be1),
	.w4(32'hbbefeb29),
	.w5(32'hbc0a5eff),
	.w6(32'h3b0e6740),
	.w7(32'h3bc3d2a7),
	.w8(32'h3b7e988e),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b74fe17),
	.w1(32'hbbada540),
	.w2(32'hbc032bc2),
	.w3(32'hbb2f8c48),
	.w4(32'h3a4c0fe5),
	.w5(32'h3b9c8051),
	.w6(32'hbc00f787),
	.w7(32'hbc432886),
	.w8(32'hbc3b87c4),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1de9fd),
	.w1(32'hbc7ad15c),
	.w2(32'h37bf7692),
	.w3(32'hbb44aa2a),
	.w4(32'h3c3b1f78),
	.w5(32'h3c865ebb),
	.w6(32'h3c519942),
	.w7(32'h3cfdfa90),
	.w8(32'h3ca9c47b),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af3a5f8),
	.w1(32'h3a5a65c6),
	.w2(32'h3acb2ac0),
	.w3(32'hb9fce9b7),
	.w4(32'h39c38a7e),
	.w5(32'hba1609cf),
	.w6(32'hbb95196d),
	.w7(32'hbb55b3db),
	.w8(32'hbbbd9ace),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390440fe),
	.w1(32'hbadd4de4),
	.w2(32'hb9846775),
	.w3(32'h3b24e71b),
	.w4(32'hbb0af107),
	.w5(32'hbb063181),
	.w6(32'hba04f8b6),
	.w7(32'h3b43c2e1),
	.w8(32'h3b9e4fa4),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb716381),
	.w1(32'hbb2915de),
	.w2(32'hbbc50791),
	.w3(32'h3a5e8816),
	.w4(32'h3b9eadde),
	.w5(32'h3c17a4f6),
	.w6(32'hbbc7298d),
	.w7(32'hbb94bf41),
	.w8(32'hbc0c8f3c),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc399da),
	.w1(32'hbc71be38),
	.w2(32'hbc12b45f),
	.w3(32'h3b650f32),
	.w4(32'hbc238fd7),
	.w5(32'hbc539e14),
	.w6(32'hbb645415),
	.w7(32'h3a8d6af5),
	.w8(32'h39eddcb2),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbe4646),
	.w1(32'hbc7e6cf5),
	.w2(32'hbbaa1a0a),
	.w3(32'hbc4c2824),
	.w4(32'h3c029096),
	.w5(32'h3c3f09e6),
	.w6(32'hbc18d7a4),
	.w7(32'hbbb1e658),
	.w8(32'hbc90e3ff),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad7eee6),
	.w1(32'hbb35de84),
	.w2(32'h3b354ba2),
	.w3(32'h3be32776),
	.w4(32'h3bb20b21),
	.w5(32'h3b8e4f7b),
	.w6(32'h3ba07a6a),
	.w7(32'h3c33420f),
	.w8(32'hbb59c93f),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf3123e),
	.w1(32'hbc0c68c3),
	.w2(32'h3b0a8688),
	.w3(32'h3bb40715),
	.w4(32'hbcf7bc93),
	.w5(32'hbc8ae8d6),
	.w6(32'h3b4ef531),
	.w7(32'h3cfcc6b1),
	.w8(32'h3d4ecbee),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c093da6),
	.w1(32'h3c43dc83),
	.w2(32'h3b195ea0),
	.w3(32'hbbd20434),
	.w4(32'h3c5238fa),
	.w5(32'h3bee6766),
	.w6(32'h3bf4d23f),
	.w7(32'h3b110c83),
	.w8(32'h38ebf3b9),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb251ee1),
	.w1(32'h3b2fc5e6),
	.w2(32'h3ba19a1d),
	.w3(32'hba208292),
	.w4(32'h3af71970),
	.w5(32'h3b7653ef),
	.w6(32'hbb584246),
	.w7(32'hbbcf1993),
	.w8(32'hbbd6cb8a),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb037867),
	.w1(32'hbb215fa0),
	.w2(32'h3b9b2b2a),
	.w3(32'h39baa151),
	.w4(32'hbbe32d99),
	.w5(32'h39accd64),
	.w6(32'hbaab2682),
	.w7(32'hbad69985),
	.w8(32'hbab98a4c),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc892d45),
	.w1(32'hbbe6771f),
	.w2(32'h3b8a0c6e),
	.w3(32'hbb208abb),
	.w4(32'h3b8f5d3f),
	.w5(32'hbba619c3),
	.w6(32'h3bf0b860),
	.w7(32'h3c2b3dc2),
	.w8(32'h3b147164),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8c6727),
	.w1(32'h3b2f0705),
	.w2(32'h3bb1f230),
	.w3(32'hbb3f88d0),
	.w4(32'hbba6e9a6),
	.w5(32'hbbde4c57),
	.w6(32'h3b8d26ac),
	.w7(32'h380a8551),
	.w8(32'h3b819792),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b302923),
	.w1(32'h39f45a9d),
	.w2(32'h38fb8863),
	.w3(32'hbbbe392b),
	.w4(32'hbca34823),
	.w5(32'hbc9c9e59),
	.w6(32'h3c8851f5),
	.w7(32'h3ca11c7b),
	.w8(32'h3c96d576),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b942b4c),
	.w1(32'hb6c18582),
	.w2(32'h3b357346),
	.w3(32'hbc6b8932),
	.w4(32'hba4fedfd),
	.w5(32'hbb234209),
	.w6(32'h3ba8c85e),
	.w7(32'h3aaeb391),
	.w8(32'h3b47fda8),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9d2b36),
	.w1(32'hbbfc283b),
	.w2(32'hb9a89ec4),
	.w3(32'hbbb461c2),
	.w4(32'hbac97e78),
	.w5(32'h3ab152b2),
	.w6(32'h3c4670d6),
	.w7(32'h3cb9d895),
	.w8(32'h3ca80cc2),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9cc7bc),
	.w1(32'hbc444883),
	.w2(32'hbbb0a941),
	.w3(32'hbc6db6d5),
	.w4(32'hba513d98),
	.w5(32'h3c014cd0),
	.w6(32'hbc260d37),
	.w7(32'hbbfcc416),
	.w8(32'h3bb242f6),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9a9f4b),
	.w1(32'hbbdf408c),
	.w2(32'hbbb880dc),
	.w3(32'hbb55c855),
	.w4(32'hbc152a6f),
	.w5(32'hbb583be3),
	.w6(32'hbb7b0983),
	.w7(32'hbb50a576),
	.w8(32'hbba9e94b),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba554106),
	.w1(32'h39caf09e),
	.w2(32'h3bbf6dd2),
	.w3(32'hb766de16),
	.w4(32'hbb99aae0),
	.w5(32'hbc3439d8),
	.w6(32'h3c2ed280),
	.w7(32'h3c68043d),
	.w8(32'h3c5795b7),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5e22fa),
	.w1(32'h3c735b1d),
	.w2(32'h3c7c412f),
	.w3(32'hbc5fd1fc),
	.w4(32'hbbb88ede),
	.w5(32'hbc38055b),
	.w6(32'hbb88433e),
	.w7(32'h3833e520),
	.w8(32'h39882a68),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2bccf6),
	.w1(32'hbc5fc49b),
	.w2(32'hba9363d6),
	.w3(32'hb9398053),
	.w4(32'hbcda7d90),
	.w5(32'hbc70fc9b),
	.w6(32'h3c454a6d),
	.w7(32'h3cbee94a),
	.w8(32'h3cb9c351),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd002720),
	.w1(32'hbcf305f1),
	.w2(32'hbcacece5),
	.w3(32'hbcbe8535),
	.w4(32'hbba24ae9),
	.w5(32'hbc985cd8),
	.w6(32'h3bb5f308),
	.w7(32'h3d1b9608),
	.w8(32'h3bd0cefe),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd25294c),
	.w1(32'hbca957c9),
	.w2(32'hbb212392),
	.w3(32'hbc8d8a3e),
	.w4(32'hbc62264e),
	.w5(32'hbbee5aee),
	.w6(32'h3c4477c9),
	.w7(32'h3d055911),
	.w8(32'h3ce5213a),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb512eb9),
	.w1(32'hbc5628e4),
	.w2(32'hbbf9480f),
	.w3(32'hbccc74db),
	.w4(32'hbc84c7e2),
	.w5(32'hbc179971),
	.w6(32'hbb476a65),
	.w7(32'hbae71703),
	.w8(32'h3c3357d7),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcafb7a2),
	.w1(32'h3beaea4e),
	.w2(32'h3b03431a),
	.w3(32'hbc8a3d5f),
	.w4(32'h3b0c09fd),
	.w5(32'h3a7276a7),
	.w6(32'h3990b027),
	.w7(32'hbb360678),
	.w8(32'h39fca55b),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a86a20f),
	.w1(32'hbb03542c),
	.w2(32'hbbac4d01),
	.w3(32'h3a1f26f2),
	.w4(32'h3a461185),
	.w5(32'hbb01a52b),
	.w6(32'h3baf0dcd),
	.w7(32'h3bb0b971),
	.w8(32'h3b52fa1b),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e2a409),
	.w1(32'h3b84d971),
	.w2(32'h3ba352db),
	.w3(32'hba82cdca),
	.w4(32'h3bbca091),
	.w5(32'h3c17a6c1),
	.w6(32'hbbae599f),
	.w7(32'hbb72f248),
	.w8(32'hb991207c),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6d6542),
	.w1(32'h3aef32c0),
	.w2(32'h3c0c983c),
	.w3(32'h3c2edac3),
	.w4(32'hbbc83f61),
	.w5(32'hbbf07639),
	.w6(32'h3b68fccd),
	.w7(32'h3c179770),
	.w8(32'h3c39f288),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c01c6b9),
	.w1(32'hbb84581c),
	.w2(32'h39c9a8ec),
	.w3(32'hbafcd3df),
	.w4(32'hbb24af21),
	.w5(32'h3c0402a2),
	.w6(32'hbb947ff7),
	.w7(32'hbbdc61ff),
	.w8(32'hbc17fccf),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbad39e5),
	.w1(32'hbb844502),
	.w2(32'hbbb28845),
	.w3(32'hbb4fa76a),
	.w4(32'h3c1497a3),
	.w5(32'h3c776214),
	.w6(32'hbb9bbeec),
	.w7(32'hbc54c38b),
	.w8(32'hbc552dd7),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3822a461),
	.w1(32'h3c5162a6),
	.w2(32'h3b2aebac),
	.w3(32'h3ae3a3c8),
	.w4(32'hbb95eced),
	.w5(32'hbc230753),
	.w6(32'h37b20452),
	.w7(32'h3b2541d1),
	.w8(32'hbb54190e),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbba5e6e),
	.w1(32'hbb83dd87),
	.w2(32'h3a5b003a),
	.w3(32'hba906043),
	.w4(32'h3ad72126),
	.w5(32'h3bdea910),
	.w6(32'hbadf7f48),
	.w7(32'h3abe2791),
	.w8(32'hb856c557),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e2914),
	.w1(32'hba86b031),
	.w2(32'hbb80148b),
	.w3(32'h3ba28fd9),
	.w4(32'hbb9e6704),
	.w5(32'hbc542ee4),
	.w6(32'hbb851ed7),
	.w7(32'h3b6ba3f9),
	.w8(32'h3c089b3b),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb024a46),
	.w1(32'hbc719678),
	.w2(32'hbb41cb98),
	.w3(32'hbbd6c162),
	.w4(32'hbc76d275),
	.w5(32'hbb81322c),
	.w6(32'hbb4e86b0),
	.w7(32'h3b125ce2),
	.w8(32'h3bad0899),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb41e573),
	.w1(32'h3a3acd6d),
	.w2(32'h3b676166),
	.w3(32'h3a1fd476),
	.w4(32'hbbd796fc),
	.w5(32'hbc3c1a61),
	.w6(32'h3c31cf8a),
	.w7(32'h3cefa088),
	.w8(32'h3c3f985a),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4afd9f),
	.w1(32'hbad9b1c7),
	.w2(32'hb9eebdd2),
	.w3(32'h3ace0364),
	.w4(32'hbbc46fa2),
	.w5(32'hbc00f10b),
	.w6(32'h3b6b0e33),
	.w7(32'h3bba0950),
	.w8(32'hb9c60e04),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba722efc),
	.w1(32'hbb5760b7),
	.w2(32'h3a18df60),
	.w3(32'hbb90f6b2),
	.w4(32'hbb14fb6b),
	.w5(32'h3b7cf8f5),
	.w6(32'hbb6305a8),
	.w7(32'hbbaecb3e),
	.w8(32'hbbb6753d),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc0bd43),
	.w1(32'h3b9398da),
	.w2(32'hbb00f1fb),
	.w3(32'hbb027945),
	.w4(32'hbc848902),
	.w5(32'hbb960336),
	.w6(32'hbae3b726),
	.w7(32'h3ad4db7d),
	.w8(32'hbb6348c9),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadaa754),
	.w1(32'hbbefa7f5),
	.w2(32'hbc5fe4c7),
	.w3(32'hbb9381d8),
	.w4(32'hbc85052a),
	.w5(32'hbc4b48a4),
	.w6(32'hbb72af5f),
	.w7(32'hbb9b0d21),
	.w8(32'hbc189649),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0339f8),
	.w1(32'h3b04dc8e),
	.w2(32'h3b71d8c4),
	.w3(32'hbb8ca6bb),
	.w4(32'hbc1dc9c9),
	.w5(32'hbc880511),
	.w6(32'h3bad08ab),
	.w7(32'h3ca738e2),
	.w8(32'h3c81ed1a),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7e87ac),
	.w1(32'h3ac4822b),
	.w2(32'h3c25be5a),
	.w3(32'hbbd338b8),
	.w4(32'h3b4fdad4),
	.w5(32'h3b91873c),
	.w6(32'hbb7616b0),
	.w7(32'hbb9b162b),
	.w8(32'hbba4295a),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba5c0d3),
	.w1(32'h3c6f18d5),
	.w2(32'h3b8709a5),
	.w3(32'hbaf7d13d),
	.w4(32'hbc103ecb),
	.w5(32'hbc39c6e8),
	.w6(32'hbbcc93f6),
	.w7(32'hbb58989a),
	.w8(32'hbbd78a25),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c280554),
	.w1(32'hbad2e7a9),
	.w2(32'hbb401c78),
	.w3(32'hba0d4aac),
	.w4(32'hbc22f383),
	.w5(32'hbc20cbba),
	.w6(32'hbc006b65),
	.w7(32'hbb5652c8),
	.w8(32'hbb009d2f),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc232103),
	.w1(32'hbc496818),
	.w2(32'hbb1ad485),
	.w3(32'hbc21f92e),
	.w4(32'hbc1e07ff),
	.w5(32'h390634b6),
	.w6(32'hbb628e53),
	.w7(32'h3bd87cca),
	.w8(32'h3c435ece),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a06176e),
	.w1(32'hbb01639e),
	.w2(32'h3aae2fc2),
	.w3(32'h3ad5ed67),
	.w4(32'hbb5f9e19),
	.w5(32'h3b0ac1c2),
	.w6(32'h3a2bdd38),
	.w7(32'h39c15833),
	.w8(32'h3b657dc4),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf837ea),
	.w1(32'h3bef3c66),
	.w2(32'hbba95447),
	.w3(32'h3b9c714a),
	.w4(32'hbbbd7807),
	.w5(32'hbc077f1b),
	.w6(32'hbb6c6378),
	.w7(32'hbba37df0),
	.w8(32'hbb807fc9),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0ec967),
	.w1(32'h3bce826f),
	.w2(32'h3b08409a),
	.w3(32'hbbf6b4ef),
	.w4(32'h3cb6517c),
	.w5(32'h3d00dff5),
	.w6(32'hbbfe0f28),
	.w7(32'hbca0358c),
	.w8(32'hbc9367bf),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0b67b6),
	.w1(32'hba8cee30),
	.w2(32'hba498ef8),
	.w3(32'h3c9f03b0),
	.w4(32'h39fcf0c1),
	.w5(32'h3b05055e),
	.w6(32'hbb73a5c0),
	.w7(32'hbb351b0e),
	.w8(32'hbaa339ef),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba87f884),
	.w1(32'hb9cd5319),
	.w2(32'hbbc432a7),
	.w3(32'h3b984d0a),
	.w4(32'h395f0ca0),
	.w5(32'h3b40d03a),
	.w6(32'hbb58daf8),
	.w7(32'hbbb1e6e1),
	.w8(32'hbc4576f3),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca1aa26),
	.w1(32'hbb3c80c9),
	.w2(32'hbb96a221),
	.w3(32'hb9b908d7),
	.w4(32'hbaaee618),
	.w5(32'hbb404103),
	.w6(32'hbb9038d5),
	.w7(32'hbb40ce02),
	.w8(32'hbbf21e3a),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98601c3),
	.w1(32'h3b881e9e),
	.w2(32'h3c016b80),
	.w3(32'hbb135cd9),
	.w4(32'hbb968da7),
	.w5(32'h3ad21cf6),
	.w6(32'hbb8f2b1a),
	.w7(32'hba03388d),
	.w8(32'h3ae49f5f),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6dc7f6),
	.w1(32'h3b90cfd0),
	.w2(32'h3bfcd0a6),
	.w3(32'h3b9ca498),
	.w4(32'hbb06876d),
	.w5(32'hba50b0de),
	.w6(32'h3b484062),
	.w7(32'h3a3505b1),
	.w8(32'h3b4551a3),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2a8271),
	.w1(32'h3ba5e191),
	.w2(32'h3b5fa96e),
	.w3(32'h3a859bf3),
	.w4(32'h3bed5e34),
	.w5(32'h3c311b01),
	.w6(32'h38f55269),
	.w7(32'hb93ed095),
	.w8(32'hba0f9267),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1fcb31),
	.w1(32'hba35c662),
	.w2(32'h39e36184),
	.w3(32'h3b92a683),
	.w4(32'hba5f761b),
	.w5(32'hba2e5f4a),
	.w6(32'h3504cc7d),
	.w7(32'h3b3789ed),
	.w8(32'h3ba701ad),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6fae54),
	.w1(32'h3ba259f0),
	.w2(32'h3baa9e84),
	.w3(32'h3ac57959),
	.w4(32'hbba0fed1),
	.w5(32'hbb9f742e),
	.w6(32'h3c005d4c),
	.w7(32'h3c03a7a3),
	.w8(32'h3c546448),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fe0645),
	.w1(32'hbbeeda89),
	.w2(32'h3a0c4993),
	.w3(32'hbb1d1ee3),
	.w4(32'hbbd5c6f4),
	.w5(32'h3b210922),
	.w6(32'h3ba330e3),
	.w7(32'h3c75034c),
	.w8(32'h3c1e0413),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba8c093),
	.w1(32'h39834d36),
	.w2(32'h3ab1c9d5),
	.w3(32'h3a10f54a),
	.w4(32'hbbc5cda0),
	.w5(32'hbc27aac2),
	.w6(32'h38de2cc0),
	.w7(32'h3c50abc6),
	.w8(32'h3b72b05b),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3421ce),
	.w1(32'hba08782e),
	.w2(32'hba3f6989),
	.w3(32'hbc86dc61),
	.w4(32'hba450ae2),
	.w5(32'hb8d15460),
	.w6(32'h3a838c8b),
	.w7(32'hbad59834),
	.w8(32'hbb00678c),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa8f15e),
	.w1(32'h3c39abfc),
	.w2(32'h3c51f73a),
	.w3(32'hbc6034e3),
	.w4(32'hbad349f7),
	.w5(32'hbb5c30ab),
	.w6(32'hb9df34ec),
	.w7(32'h39741644),
	.w8(32'h3bea1300),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0559d3),
	.w1(32'h3b0f0b75),
	.w2(32'h3be50433),
	.w3(32'h3c0a7c2c),
	.w4(32'h3b878ae7),
	.w5(32'h3bde2ae3),
	.w6(32'h3bbd6eea),
	.w7(32'h3bdb76ec),
	.w8(32'h39f59ad1),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8a60f9),
	.w1(32'h3b263546),
	.w2(32'h3a41d187),
	.w3(32'hbbb0ed21),
	.w4(32'h3b37a0eb),
	.w5(32'h3bc42a59),
	.w6(32'hbb4cbed8),
	.w7(32'hbb701bfb),
	.w8(32'hbc0e52b5),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8856e8),
	.w1(32'h3b3d7c19),
	.w2(32'h3bd79dcc),
	.w3(32'h3ba99310),
	.w4(32'hbb4c2d04),
	.w5(32'h3b130486),
	.w6(32'h3a0bb142),
	.w7(32'h3c0bd5d2),
	.w8(32'h3ba92349),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b83eb5a),
	.w1(32'h3bd69d59),
	.w2(32'h3c0f17ae),
	.w3(32'hbade1814),
	.w4(32'h3bf67fc0),
	.w5(32'h3b272330),
	.w6(32'h3bf4f77e),
	.w7(32'h3c0ce7aa),
	.w8(32'h39f963ab),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba42f1a),
	.w1(32'hbbc9c1b6),
	.w2(32'hbbd01f55),
	.w3(32'h3a523252),
	.w4(32'hbc323aa2),
	.w5(32'hbbb3065e),
	.w6(32'hbae5bab2),
	.w7(32'h3aa4b4c3),
	.w8(32'h3ab64e74),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1cfa26),
	.w1(32'hbb56b065),
	.w2(32'hb9281237),
	.w3(32'hbb51cbab),
	.w4(32'hba8cd67b),
	.w5(32'hbb0ee7d6),
	.w6(32'hbb3d5373),
	.w7(32'hbb279ea5),
	.w8(32'hbafd45d1),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae807ab),
	.w1(32'h3aafde19),
	.w2(32'hbc139a79),
	.w3(32'hbb74eba7),
	.w4(32'hbb7d0ed5),
	.w5(32'hbb33e477),
	.w6(32'hbae08036),
	.w7(32'hbb6fa749),
	.w8(32'h3ac0f5b1),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule