module layer_8_featuremap_215(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b40011a),
	.w1(32'hbbbc1564),
	.w2(32'hbb4bdd9e),
	.w3(32'h3bac1d08),
	.w4(32'hbb57ddf2),
	.w5(32'h3bc39d3c),
	.w6(32'h3c3e5268),
	.w7(32'h3b48adc4),
	.w8(32'h3b7f9e38),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1b1db8),
	.w1(32'hbb665500),
	.w2(32'h3b186932),
	.w3(32'hbb9a84a5),
	.w4(32'hbb450fe4),
	.w5(32'h3aef8b7c),
	.w6(32'hbb47a519),
	.w7(32'hbb17f431),
	.w8(32'hba95ecce),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b087ab4),
	.w1(32'h368e1090),
	.w2(32'hbc7f45ed),
	.w3(32'h3a85b9a6),
	.w4(32'h3c2715bf),
	.w5(32'hbc020278),
	.w6(32'h37835637),
	.w7(32'hbbe5e7ca),
	.w8(32'hbbf7e460),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf04f08),
	.w1(32'h3bae04e7),
	.w2(32'hbbde1e17),
	.w3(32'hbc60e14c),
	.w4(32'h3b8c3c4c),
	.w5(32'hbc98e5e0),
	.w6(32'hbc397ac2),
	.w7(32'h3b71796b),
	.w8(32'h3ad29f46),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6774f5),
	.w1(32'hb9f606ee),
	.w2(32'h3b465733),
	.w3(32'h3b05c244),
	.w4(32'hbad11224),
	.w5(32'h3b1ee526),
	.w6(32'h3abfc756),
	.w7(32'h3b8e01de),
	.w8(32'h3ade6eec),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af8eb57),
	.w1(32'h3ba820aa),
	.w2(32'h3cc76f45),
	.w3(32'h3a56a2a9),
	.w4(32'hbb350b10),
	.w5(32'h3c9eeea6),
	.w6(32'h3bec190b),
	.w7(32'hbb82cc10),
	.w8(32'hbac5db6e),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af94d60),
	.w1(32'h3b11fabd),
	.w2(32'h39cf2cd6),
	.w3(32'h3bea9355),
	.w4(32'h3a4c1a7a),
	.w5(32'hba514536),
	.w6(32'h3a23356d),
	.w7(32'h3a6f912b),
	.w8(32'h3b379b83),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b14d8d1),
	.w1(32'hbc060048),
	.w2(32'hbc6779a4),
	.w3(32'h3ba77574),
	.w4(32'h39a04f01),
	.w5(32'hbc1530fc),
	.w6(32'h3c392725),
	.w7(32'hbc5eb1d5),
	.w8(32'hb98e7af0),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4f0326),
	.w1(32'h3afac840),
	.w2(32'h3bf3115e),
	.w3(32'h3b3153d7),
	.w4(32'h3b9c859e),
	.w5(32'h3bd1f280),
	.w6(32'h39283bc7),
	.w7(32'h3a987043),
	.w8(32'hba821a6a),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba43943),
	.w1(32'h3b5cd02e),
	.w2(32'h3b06ba9e),
	.w3(32'h3b9d0ff1),
	.w4(32'h3b987ccc),
	.w5(32'hba63067e),
	.w6(32'h3aa579f4),
	.w7(32'h3b3dd6c3),
	.w8(32'hba249fc4),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39424c5e),
	.w1(32'hbbefdce9),
	.w2(32'hbbee9878),
	.w3(32'h3c25e184),
	.w4(32'hbc4e1e73),
	.w5(32'hbc7fbb84),
	.w6(32'hbc1296e3),
	.w7(32'hbbd31e70),
	.w8(32'hbbdc5fb4),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb397e3e),
	.w1(32'hbba6cf9a),
	.w2(32'hbc10610b),
	.w3(32'hbbb1186f),
	.w4(32'hbbb38c1a),
	.w5(32'h39c53db4),
	.w6(32'hbbeab567),
	.w7(32'hbba80b47),
	.w8(32'h3a907cdf),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9f5db9),
	.w1(32'hbc824179),
	.w2(32'hbc1f134c),
	.w3(32'h3b7a10bc),
	.w4(32'hbc0672b1),
	.w5(32'hbc6ed058),
	.w6(32'hbb514aae),
	.w7(32'hbb9d60fa),
	.w8(32'hbacae19e),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc17372c),
	.w1(32'h3a37f7e0),
	.w2(32'hbbc3250a),
	.w3(32'hbb9b99a9),
	.w4(32'hba9e0a6e),
	.w5(32'hbc04a34a),
	.w6(32'hbb799771),
	.w7(32'hbb673414),
	.w8(32'hbba2de84),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9cb211),
	.w1(32'hbb3a4c34),
	.w2(32'hbbd1e0bb),
	.w3(32'hbb93bd05),
	.w4(32'hba85e357),
	.w5(32'hbb6672b5),
	.w6(32'hbb513090),
	.w7(32'hbb921d38),
	.w8(32'hb9f8815d),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a81fd09),
	.w1(32'hbcde876e),
	.w2(32'h3c87f174),
	.w3(32'h3b23e8e7),
	.w4(32'hbca5cf86),
	.w5(32'h3cdced53),
	.w6(32'hbc65f0d2),
	.w7(32'h3b382011),
	.w8(32'h3b1af3f6),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb79a3c2),
	.w1(32'h3bcd88a7),
	.w2(32'hbc19d2bc),
	.w3(32'hbaadb1aa),
	.w4(32'h3cb86e3c),
	.w5(32'h3c0e04ea),
	.w6(32'h3b0f2469),
	.w7(32'h3a9454cd),
	.w8(32'h3ba45d1f),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbef317a),
	.w1(32'hbb2d829c),
	.w2(32'hbba8b74a),
	.w3(32'h3bd572ea),
	.w4(32'hba3c075d),
	.w5(32'h3b5e0892),
	.w6(32'hbb8210fa),
	.w7(32'hbaa38d45),
	.w8(32'h3b13caeb),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9780ca3),
	.w1(32'hbc497565),
	.w2(32'h3c13efb7),
	.w3(32'hbb87201b),
	.w4(32'hba4af06b),
	.w5(32'hbb7fea61),
	.w6(32'h3b6a62db),
	.w7(32'h3a9d5a24),
	.w8(32'h3c64de39),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b92465c),
	.w1(32'h3b92eac4),
	.w2(32'hbaaef02f),
	.w3(32'h3abfe8bb),
	.w4(32'h3b568043),
	.w5(32'h3a15565e),
	.w6(32'hba8a064a),
	.w7(32'hbb14a023),
	.w8(32'hba6aebe8),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0eb559),
	.w1(32'h3e034a61),
	.w2(32'hbb680686),
	.w3(32'hba487707),
	.w4(32'h3dd36d1f),
	.w5(32'h3c2a1380),
	.w6(32'h3d0450f8),
	.w7(32'hbc3c7eab),
	.w8(32'hbc4086f5),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcfca4de),
	.w1(32'hb9eabbeb),
	.w2(32'hbbe20bbd),
	.w3(32'hbcb56503),
	.w4(32'hbbe09a9c),
	.w5(32'h3c4a2b7f),
	.w6(32'h3c1831c6),
	.w7(32'hbc062550),
	.w8(32'h3aa6be11),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd92c42),
	.w1(32'hbb769b1e),
	.w2(32'hbc5732fa),
	.w3(32'hbada8397),
	.w4(32'hbad2c1b9),
	.w5(32'hbbb0e2fd),
	.w6(32'hbbf1306a),
	.w7(32'hbc4d505a),
	.w8(32'h3b00a5e4),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba9d87e),
	.w1(32'h3bcb2efa),
	.w2(32'hbbe1cab0),
	.w3(32'h3b67ed75),
	.w4(32'h3b5086e5),
	.w5(32'hbc1f73db),
	.w6(32'hba7eb282),
	.w7(32'hbb4534dc),
	.w8(32'h3b25a455),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb514629),
	.w1(32'h3bfe2206),
	.w2(32'h3ab4890f),
	.w3(32'hbc08b1cd),
	.w4(32'h3aaf659a),
	.w5(32'h3b0b4d21),
	.w6(32'h3c335104),
	.w7(32'h3ae49d88),
	.w8(32'h3aee42e3),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b280c86),
	.w1(32'h3dd057af),
	.w2(32'h3b32b8cc),
	.w3(32'hbb5ae16e),
	.w4(32'h3c569025),
	.w5(32'h3ca7d536),
	.w6(32'h3d895835),
	.w7(32'hbc8f227d),
	.w8(32'hbc998e1c),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcec8f21),
	.w1(32'h3c2fddba),
	.w2(32'h3c0a55aa),
	.w3(32'hbc2580d4),
	.w4(32'h3c447027),
	.w5(32'h3c0bdfe3),
	.w6(32'h3bfa0375),
	.w7(32'h3a7e1bea),
	.w8(32'h3b9b8950),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2c68ad),
	.w1(32'h3c3e0ccc),
	.w2(32'hbca90657),
	.w3(32'hbc43c3e1),
	.w4(32'h3caa9f41),
	.w5(32'hbc01926b),
	.w6(32'hbc01cf39),
	.w7(32'hbbbf3f18),
	.w8(32'hbc08cfdb),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbafbcfa),
	.w1(32'h3bfb8b41),
	.w2(32'hbb7ad51f),
	.w3(32'hbbace09d),
	.w4(32'h3be1a4a1),
	.w5(32'h391dc6d0),
	.w6(32'h3bc2140a),
	.w7(32'hbc1c6b0b),
	.w8(32'hbb80a4b9),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b7ba2),
	.w1(32'hbb6870d6),
	.w2(32'hbbea2c71),
	.w3(32'hbb4cdf9e),
	.w4(32'hbb70569c),
	.w5(32'hbbce1144),
	.w6(32'h399e8ad0),
	.w7(32'hbb1c8460),
	.w8(32'h3bd89e40),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba1bd9a),
	.w1(32'h3c263a21),
	.w2(32'h3ae5b421),
	.w3(32'h3bcabce9),
	.w4(32'h3b7c0477),
	.w5(32'hbb209f4d),
	.w6(32'h3bc85cd8),
	.w7(32'h3b81acb6),
	.w8(32'hbb170a1c),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6c68fe),
	.w1(32'h3cc05889),
	.w2(32'hbb00b652),
	.w3(32'h3b431b7a),
	.w4(32'h3c86f8c7),
	.w5(32'h3b9338ce),
	.w6(32'hbaa940b9),
	.w7(32'hbc380b9c),
	.w8(32'hbcb14011),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcab147c),
	.w1(32'hba1f0caa),
	.w2(32'h3b00fdc5),
	.w3(32'hbc949ac2),
	.w4(32'h3bc26cfd),
	.w5(32'hbab3a757),
	.w6(32'hbb20a058),
	.w7(32'h3bdfcfaa),
	.w8(32'h3bc0d2b5),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c21e5c0),
	.w1(32'h3af6cd8c),
	.w2(32'hbb7f3290),
	.w3(32'h3b5e9826),
	.w4(32'h3bbd5d20),
	.w5(32'hba9b6d2b),
	.w6(32'h3ad94463),
	.w7(32'h3b174ffd),
	.w8(32'h3739b9a2),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39275463),
	.w1(32'hbbad18fb),
	.w2(32'hbbd47c05),
	.w3(32'hb8890f00),
	.w4(32'hb9d02378),
	.w5(32'h3a91e0d9),
	.w6(32'hbaec02fd),
	.w7(32'hbb282441),
	.w8(32'h3a93b9e7),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398ec3f1),
	.w1(32'h3c262db3),
	.w2(32'hbc31df06),
	.w3(32'h3b2204ea),
	.w4(32'h3c0c2440),
	.w5(32'hbb21f678),
	.w6(32'h3b58c4af),
	.w7(32'hbaa72d4a),
	.w8(32'hba8837ab),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39773744),
	.w1(32'h39d0e3ec),
	.w2(32'h3bde690a),
	.w3(32'hbb581390),
	.w4(32'h3b027da6),
	.w5(32'h3ba39234),
	.w6(32'h3b290541),
	.w7(32'h3b947b92),
	.w8(32'h3baf3cf2),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c09d506),
	.w1(32'hbb31928f),
	.w2(32'h3b196992),
	.w3(32'h3c043b5f),
	.w4(32'h3b4236c9),
	.w5(32'h3bb9ad12),
	.w6(32'h3a966f9e),
	.w7(32'h3b5451ee),
	.w8(32'h3b2ab003),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba934cf),
	.w1(32'hbabe370e),
	.w2(32'hba24c1c2),
	.w3(32'h3be928c3),
	.w4(32'h3bc62815),
	.w5(32'h3c2590e7),
	.w6(32'hbb75aab4),
	.w7(32'hbb862b49),
	.w8(32'h3941e035),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b24b27a),
	.w1(32'h3b0ecad0),
	.w2(32'hbbdbab61),
	.w3(32'h3ac45e8b),
	.w4(32'hbab3da6a),
	.w5(32'hbbdf28e7),
	.w6(32'h3b91482c),
	.w7(32'hbb43c6ad),
	.w8(32'h3add1742),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba6c382),
	.w1(32'h3b024e8c),
	.w2(32'h3b8a7a7c),
	.w3(32'hbc1243af),
	.w4(32'h3bbf0bce),
	.w5(32'h3bf62c5b),
	.w6(32'h39af2ab3),
	.w7(32'h3afa55a6),
	.w8(32'h3b4b5459),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba2a3e1),
	.w1(32'hbc00b78b),
	.w2(32'h3bdcc53c),
	.w3(32'h3bdf6f3e),
	.w4(32'hbb988cf1),
	.w5(32'h3be18144),
	.w6(32'hbbae53de),
	.w7(32'h3be29c69),
	.w8(32'h3b653330),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3fb9c3),
	.w1(32'hb950beea),
	.w2(32'h3bc282f1),
	.w3(32'h3b96c7cf),
	.w4(32'h3a8bcc8a),
	.w5(32'h3bfd3db8),
	.w6(32'h3b856029),
	.w7(32'h3b25c0dd),
	.w8(32'hbbd4e6d0),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad490cb),
	.w1(32'hbc434f63),
	.w2(32'h3ae18ccf),
	.w3(32'hbacce9df),
	.w4(32'hbc4c4f3b),
	.w5(32'hba91c8c8),
	.w6(32'hbc3805f1),
	.w7(32'hb91ebe89),
	.w8(32'hbb978dc2),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb127204),
	.w1(32'hbbdd94d0),
	.w2(32'hbc8c58ab),
	.w3(32'h3bb8054a),
	.w4(32'hbb4a6eff),
	.w5(32'hbcb187b7),
	.w6(32'hbc1e9202),
	.w7(32'hbc083bf0),
	.w8(32'h3bb248e0),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1c4d16),
	.w1(32'h37e2bc37),
	.w2(32'hbb1bcc4a),
	.w3(32'h3ba030f5),
	.w4(32'h3b925673),
	.w5(32'h3b15b363),
	.w6(32'hbb2f8d34),
	.w7(32'hbb565743),
	.w8(32'h3a76f56c),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba1e75c),
	.w1(32'hbc4513bc),
	.w2(32'hbc4cc2a1),
	.w3(32'h3bcaa334),
	.w4(32'hbc8abe4e),
	.w5(32'hbc7ccf56),
	.w6(32'hbc3c13bd),
	.w7(32'hbc2c99e0),
	.w8(32'hbc0f6dd6),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba80314),
	.w1(32'h3be56da0),
	.w2(32'hbc365826),
	.w3(32'hbc26c196),
	.w4(32'h3ac09d87),
	.w5(32'hb9128987),
	.w6(32'h3b4a0401),
	.w7(32'hbb35f528),
	.w8(32'h3a674e98),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbfbf5b),
	.w1(32'h3c0ebc64),
	.w2(32'hbc12cba9),
	.w3(32'hbb8848ab),
	.w4(32'h3c2e468f),
	.w5(32'h3bd79100),
	.w6(32'h3c3a6079),
	.w7(32'hbc05aba8),
	.w8(32'h3b982618),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa284eb),
	.w1(32'h3c886289),
	.w2(32'h3c93802f),
	.w3(32'hba9eb873),
	.w4(32'h3cb2f402),
	.w5(32'h3c77058b),
	.w6(32'h3c3c16d0),
	.w7(32'hbae200d3),
	.w8(32'hbb23005b),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc572816),
	.w1(32'hbb6e8587),
	.w2(32'hbb07b2c1),
	.w3(32'hbbe2a593),
	.w4(32'hbbc3306c),
	.w5(32'hbb9bbd93),
	.w6(32'hbb8348a7),
	.w7(32'hbb5d5e63),
	.w8(32'hbb943868),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3ee0c9),
	.w1(32'hbc0c2dd7),
	.w2(32'hbb982488),
	.w3(32'h38c8e469),
	.w4(32'hbb96d1fc),
	.w5(32'hbb1bed2c),
	.w6(32'hb9aaf33c),
	.w7(32'hbaf8fbef),
	.w8(32'h3af1c071),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb01ee9),
	.w1(32'hbbdff0ca),
	.w2(32'hbb2c19b5),
	.w3(32'h3afd3cd0),
	.w4(32'hbbc2f2a9),
	.w5(32'hba8cb10d),
	.w6(32'hbae89ddd),
	.w7(32'hba897cae),
	.w8(32'hba28860e),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b02d887),
	.w1(32'h3c7b18f0),
	.w2(32'hbb5af5c0),
	.w3(32'h3ab64fe6),
	.w4(32'h3cd52924),
	.w5(32'h3a9c196f),
	.w6(32'h3c13fe8a),
	.w7(32'h3bcbf0ef),
	.w8(32'h3c45b017),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca342fe),
	.w1(32'h3b44ec98),
	.w2(32'h3c3161f3),
	.w3(32'h3c810b3a),
	.w4(32'hba71507f),
	.w5(32'h3bd4e54e),
	.w6(32'h3b81de33),
	.w7(32'h3998c95a),
	.w8(32'hbbe1894e),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb381eaa),
	.w1(32'hbbcb2512),
	.w2(32'hbbd2693f),
	.w3(32'hbb9d644e),
	.w4(32'h3b75859d),
	.w5(32'hb9c0264b),
	.w6(32'hbc76e22e),
	.w7(32'h3b301af8),
	.w8(32'hbc40873c),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4d7953),
	.w1(32'hbbeb922a),
	.w2(32'hbc01c1b8),
	.w3(32'hba8d6584),
	.w4(32'hbb2773c1),
	.w5(32'h3bbe7173),
	.w6(32'hbc5ccde8),
	.w7(32'hbc24ccfd),
	.w8(32'h3b09f706),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5dfabd),
	.w1(32'hbb87d6b4),
	.w2(32'hb9de1107),
	.w3(32'h3c504187),
	.w4(32'h3a4a4218),
	.w5(32'h3a1915eb),
	.w6(32'hbb5425db),
	.w7(32'hbab34659),
	.w8(32'h39e8bd56),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6fb562),
	.w1(32'hbb237ddc),
	.w2(32'hbbc11ee0),
	.w3(32'h3a8490bb),
	.w4(32'hbaeb72ed),
	.w5(32'hbb4076ae),
	.w6(32'hbaf1d89c),
	.w7(32'hbb43808b),
	.w8(32'h3b0639d7),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba65f4f1),
	.w1(32'hbab31fd4),
	.w2(32'hbbeffe44),
	.w3(32'h3a908b93),
	.w4(32'hbc20e59d),
	.w5(32'h3a84c286),
	.w6(32'hbbc1af88),
	.w7(32'hbb146659),
	.w8(32'h3ac65fcc),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb88e1ec),
	.w1(32'hbcd2c650),
	.w2(32'hbc8dc4c4),
	.w3(32'hbb63fd5e),
	.w4(32'hbbd12a47),
	.w5(32'hba11ef1c),
	.w6(32'hbbb59250),
	.w7(32'hbc79e027),
	.w8(32'hbb412520),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb519042),
	.w1(32'h3bf3385f),
	.w2(32'h39e3cda4),
	.w3(32'hbb993faf),
	.w4(32'h3c959ca0),
	.w5(32'h3bcca373),
	.w6(32'hba7c283e),
	.w7(32'h39d1847b),
	.w8(32'hbba27520),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1f30b7),
	.w1(32'h3c648d7b),
	.w2(32'h3c39c32c),
	.w3(32'hbc072c94),
	.w4(32'h3c6cf160),
	.w5(32'h3c02aa7b),
	.w6(32'h3bd4377b),
	.w7(32'h3a10b4df),
	.w8(32'h3a46265a),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb004283),
	.w1(32'hbba33b24),
	.w2(32'hbbe619f1),
	.w3(32'h3ab73a20),
	.w4(32'hbb43eef8),
	.w5(32'hbb6091aa),
	.w6(32'hbbe30e19),
	.w7(32'hbbc5ef36),
	.w8(32'hbb5f4320),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d1779),
	.w1(32'h3b5a56cd),
	.w2(32'h3a5d1c90),
	.w3(32'hbb7e8e38),
	.w4(32'h3b2e551e),
	.w5(32'h3aebc850),
	.w6(32'h3a44b12a),
	.w7(32'hbb2495df),
	.w8(32'hba5c7887),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b03117f),
	.w1(32'hbb14594d),
	.w2(32'hbc7563db),
	.w3(32'h3b04ee98),
	.w4(32'h39fc0cfa),
	.w5(32'hbc0cb6ac),
	.w6(32'hb89bdcaa),
	.w7(32'hbba9c7cd),
	.w8(32'h3b58afdd),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb08e242),
	.w1(32'h3d120e66),
	.w2(32'hbaa277e7),
	.w3(32'hbb90877b),
	.w4(32'h3c8dcbaf),
	.w5(32'h3c310cfc),
	.w6(32'h3b186544),
	.w7(32'h3c1a985d),
	.w8(32'hbade9e7d),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6756d1),
	.w1(32'h3d407e44),
	.w2(32'hbc4b9805),
	.w3(32'hbc762e20),
	.w4(32'h3d17ec3e),
	.w5(32'h3c18f0b2),
	.w6(32'h3c9d8230),
	.w7(32'hbc5853d9),
	.w8(32'hbbb5ade9),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc241b72),
	.w1(32'hbb2b48d7),
	.w2(32'hbbdc5cac),
	.w3(32'hbc5c80be),
	.w4(32'hbad4babf),
	.w5(32'hbc217894),
	.w6(32'h3b930bd9),
	.w7(32'hbb6f55c0),
	.w8(32'hbbd4813c),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbecbf3b),
	.w1(32'h3c54a429),
	.w2(32'hbc3c4411),
	.w3(32'hbc7a2774),
	.w4(32'h3c16b184),
	.w5(32'hba4c4f23),
	.w6(32'hbae43427),
	.w7(32'hbc676991),
	.w8(32'h3b8ad952),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0d92b4),
	.w1(32'h3b06a1db),
	.w2(32'h3c99cc14),
	.w3(32'hbba0be1b),
	.w4(32'h3ba76919),
	.w5(32'h3c75355f),
	.w6(32'h3b3010b6),
	.w7(32'h3be2c2d9),
	.w8(32'hbc545246),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2f06c8),
	.w1(32'h3c6ed69e),
	.w2(32'hbad0d0e9),
	.w3(32'hbc46ebd0),
	.w4(32'h3c264ab7),
	.w5(32'hbb3840dd),
	.w6(32'h3c37a5cb),
	.w7(32'hbb140bcf),
	.w8(32'hbaa09c7b),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab30f38),
	.w1(32'h3b6f9fa0),
	.w2(32'hbc02631b),
	.w3(32'hbbe12efe),
	.w4(32'h3b2ebe52),
	.w5(32'hbbc0192e),
	.w6(32'h3c2bd45b),
	.w7(32'hbb07641b),
	.w8(32'hba8acd61),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0d83a1),
	.w1(32'h3a0d543a),
	.w2(32'hbc0a7038),
	.w3(32'hbba348fc),
	.w4(32'h3aaa542f),
	.w5(32'hbb00d773),
	.w6(32'hbc06c293),
	.w7(32'hbb78b3eb),
	.w8(32'h3afb4a3d),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be3c061),
	.w1(32'hbb504551),
	.w2(32'hbb8f394f),
	.w3(32'h3a38fb28),
	.w4(32'hbacbed5e),
	.w5(32'h3c3907f0),
	.w6(32'h3c132d1f),
	.w7(32'hbb354633),
	.w8(32'hbbd4469d),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb678273),
	.w1(32'h3a5ea6d6),
	.w2(32'h3ab8a2a0),
	.w3(32'h3abec528),
	.w4(32'h3b9e60cd),
	.w5(32'h3adcdf61),
	.w6(32'h3b9e3593),
	.w7(32'hbc480e03),
	.w8(32'hbb0671ec),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ec7421),
	.w1(32'hbabfcc8f),
	.w2(32'h3a42ed56),
	.w3(32'hba65038e),
	.w4(32'hbb38fb3e),
	.w5(32'h3be4b85b),
	.w6(32'hbb2052f2),
	.w7(32'h392da913),
	.w8(32'hb929990a),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a39812b),
	.w1(32'hbbfeb56e),
	.w2(32'h3b4d6e54),
	.w3(32'hba1a84c0),
	.w4(32'hbbeeae88),
	.w5(32'h3b8f6e29),
	.w6(32'hbb8b3391),
	.w7(32'h3b3600b4),
	.w8(32'h3b9b86b5),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8d1ee3),
	.w1(32'hbbd76a1b),
	.w2(32'hb9bc7250),
	.w3(32'h3b171c3c),
	.w4(32'h3aeeeed8),
	.w5(32'hbc4128bf),
	.w6(32'hbb34acb6),
	.w7(32'h3c078320),
	.w8(32'hbb70fafc),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba1453b),
	.w1(32'h3b8baa90),
	.w2(32'h371e6d94),
	.w3(32'hbba2e640),
	.w4(32'hbaba20e0),
	.w5(32'hbbb1ac10),
	.w6(32'h3ae3038a),
	.w7(32'hbb8422d3),
	.w8(32'hbbd3a833),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba3f0aa),
	.w1(32'h3c6a7e66),
	.w2(32'hbbb774d5),
	.w3(32'hbbb0de88),
	.w4(32'h3cc1e7d6),
	.w5(32'hbb875718),
	.w6(32'h3bd7fb09),
	.w7(32'hbbc6ca75),
	.w8(32'hbb4607d3),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc7ee89),
	.w1(32'h3c01db3a),
	.w2(32'hbb681ee2),
	.w3(32'hbc02607c),
	.w4(32'h3bd1af2c),
	.w5(32'hbb78389a),
	.w6(32'h3b70cb3a),
	.w7(32'hbb6abe5e),
	.w8(32'hbbb2c46b),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb373dec),
	.w1(32'h3bb3d7d9),
	.w2(32'hbb0cf875),
	.w3(32'hbbff68dd),
	.w4(32'h3c724436),
	.w5(32'h3c9e01ac),
	.w6(32'hbc16873e),
	.w7(32'hbc2fdb4d),
	.w8(32'h3c04b5d0),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9b65c3),
	.w1(32'hbb5ca3cb),
	.w2(32'hbc1f24a1),
	.w3(32'h3a2148bd),
	.w4(32'h3c05ab97),
	.w5(32'h3aa0d459),
	.w6(32'hbc3b7925),
	.w7(32'hbc2e48a5),
	.w8(32'hbc192772),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3d61e4),
	.w1(32'h3a7c6825),
	.w2(32'h3b242741),
	.w3(32'hbb7748bc),
	.w4(32'h3a74e4ee),
	.w5(32'hbc19c80d),
	.w6(32'hbc00faa4),
	.w7(32'h3ad2d08a),
	.w8(32'hbbb2363a),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a10e42d),
	.w1(32'h3c039689),
	.w2(32'hba099517),
	.w3(32'hba85608f),
	.w4(32'h3c3627b4),
	.w5(32'hbba474d4),
	.w6(32'hbb5ccb1d),
	.w7(32'hbbfe432a),
	.w8(32'h399ea745),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3d7d69),
	.w1(32'h3b3e1ed4),
	.w2(32'h3ba35f0c),
	.w3(32'hbc849112),
	.w4(32'h3c064900),
	.w5(32'h3b689011),
	.w6(32'h3b734af3),
	.w7(32'h3ba63379),
	.w8(32'hbb5200f1),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad3ee05),
	.w1(32'h3c1acf28),
	.w2(32'h370a0668),
	.w3(32'h3ab7d257),
	.w4(32'h3c683834),
	.w5(32'h3b6ff530),
	.w6(32'h3b2e50bb),
	.w7(32'hbb3134b4),
	.w8(32'hb850b6fc),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399fc457),
	.w1(32'hbaa21bbe),
	.w2(32'hbb4ec7cb),
	.w3(32'hbb2a63ce),
	.w4(32'h3ba70faf),
	.w5(32'h3b75521c),
	.w6(32'h3bec4839),
	.w7(32'h3b47dabf),
	.w8(32'hba9dd082),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb986b819),
	.w1(32'h3b4ab506),
	.w2(32'hbc97b0bd),
	.w3(32'h3bbb5560),
	.w4(32'hbc10433c),
	.w5(32'hbc17ad77),
	.w6(32'h3b3c9783),
	.w7(32'hbc54dd0a),
	.w8(32'h399b2353),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7cf4b1),
	.w1(32'h3c42e495),
	.w2(32'hbc023058),
	.w3(32'hbaba3be2),
	.w4(32'h3c036e4c),
	.w5(32'hbbaf14bf),
	.w6(32'h3b06754e),
	.w7(32'hbb0c73b2),
	.w8(32'hbabdd955),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6768ff),
	.w1(32'h3c248ae5),
	.w2(32'hbb7f8d18),
	.w3(32'h3b21345f),
	.w4(32'h3ae6a31b),
	.w5(32'hbb2c07ce),
	.w6(32'h3bc4e1e1),
	.w7(32'h3c2c4ead),
	.w8(32'hbad21e3a),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb306112),
	.w1(32'hbab82aeb),
	.w2(32'hba4d1866),
	.w3(32'hbbbec305),
	.w4(32'hba4e24d6),
	.w5(32'hba8f5ab7),
	.w6(32'hbb87054a),
	.w7(32'hbb44f9b2),
	.w8(32'hb94cbe4d),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb16467b),
	.w1(32'hbabf0ff3),
	.w2(32'hbb164b9d),
	.w3(32'h38c04770),
	.w4(32'hbb3a391b),
	.w5(32'hbafb1c77),
	.w6(32'hba40983d),
	.w7(32'hbb59b62b),
	.w8(32'hbb4fb9ba),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadc7418),
	.w1(32'hbc3a08f7),
	.w2(32'h3c157ea2),
	.w3(32'hbb4db622),
	.w4(32'hbc8de62b),
	.w5(32'h3c71e8bd),
	.w6(32'hbb5ed11e),
	.w7(32'hbc4b7fc3),
	.w8(32'hbbbfe3ff),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab2a689),
	.w1(32'h3a99a0bb),
	.w2(32'h3b5f13a1),
	.w3(32'h3b05b6a4),
	.w4(32'h38894721),
	.w5(32'h3bc7f009),
	.w6(32'hbb28e80c),
	.w7(32'h3727d31e),
	.w8(32'h3aaedeba),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc410e5),
	.w1(32'h3ccbbece),
	.w2(32'hbc2b868f),
	.w3(32'h3c044fc5),
	.w4(32'h3cc81aef),
	.w5(32'hbc618f48),
	.w6(32'h3b8c9441),
	.w7(32'hba2a2a83),
	.w8(32'hbbd3311f),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd2cccc),
	.w1(32'hbba1ddaf),
	.w2(32'hbb81bfae),
	.w3(32'hbc3f9651),
	.w4(32'hbba44718),
	.w5(32'hbaa878f7),
	.w6(32'hbbeb1511),
	.w7(32'hbbe5f592),
	.w8(32'hbbc091df),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbddb791),
	.w1(32'hbaf0ff81),
	.w2(32'h3b25005f),
	.w3(32'h39c875e7),
	.w4(32'h382f9e35),
	.w5(32'h3bd1f9b7),
	.w6(32'hbc51f555),
	.w7(32'hbb294bee),
	.w8(32'h3ad0d9f9),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb25e350),
	.w1(32'hbc13fc62),
	.w2(32'hbc107087),
	.w3(32'h3b65cd0f),
	.w4(32'h396e0e47),
	.w5(32'hbc2c9ac6),
	.w6(32'hbbc6f2f4),
	.w7(32'h3bdec062),
	.w8(32'h3996d438),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1cc608),
	.w1(32'h3cbc0d04),
	.w2(32'hbc4dc441),
	.w3(32'h3a7f776e),
	.w4(32'h3ca9de86),
	.w5(32'hbc67a2af),
	.w6(32'hbcb9bb5b),
	.w7(32'hba18227c),
	.w8(32'hbbdc1437),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2642d6),
	.w1(32'hbcd72757),
	.w2(32'h3c9ee5b6),
	.w3(32'h3a99abb9),
	.w4(32'hbc7a7fe7),
	.w5(32'h3c26fe92),
	.w6(32'hbbf5141c),
	.w7(32'hbba3412c),
	.w8(32'h39b2e08f),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c08f52f),
	.w1(32'h3bc6d295),
	.w2(32'h3bd102a4),
	.w3(32'h3c0081f8),
	.w4(32'h3bd7eb1e),
	.w5(32'hbbe559d8),
	.w6(32'hbb91be32),
	.w7(32'hbadf9a83),
	.w8(32'hbadb105e),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2563d5),
	.w1(32'hba21a072),
	.w2(32'hbc92d46f),
	.w3(32'h3a14dc3d),
	.w4(32'h3c376e71),
	.w5(32'hbae43a8d),
	.w6(32'hbc8e88b5),
	.w7(32'hbc9b5f35),
	.w8(32'h3a9daaa7),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4270bc),
	.w1(32'hbcaa39aa),
	.w2(32'hbbeb1412),
	.w3(32'hba206c77),
	.w4(32'hbc521a77),
	.w5(32'hb9522b92),
	.w6(32'hbcc847ef),
	.w7(32'hbbb1696a),
	.w8(32'hbbe57b88),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399c5006),
	.w1(32'h3b6a29aa),
	.w2(32'hba89bad8),
	.w3(32'hbb8efe9d),
	.w4(32'h3b7f8fd8),
	.w5(32'hb85fd98c),
	.w6(32'hbb9ba013),
	.w7(32'hbbbd13ec),
	.w8(32'hbb349a00),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f732af),
	.w1(32'h3aa66cea),
	.w2(32'h3ab1a736),
	.w3(32'h3aeeaa05),
	.w4(32'h3a9d843e),
	.w5(32'h3b773666),
	.w6(32'h3b7be8eb),
	.w7(32'h39dacd98),
	.w8(32'hbb930fa1),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4493b1),
	.w1(32'hbb902b14),
	.w2(32'h3a3e985d),
	.w3(32'h3c02e98e),
	.w4(32'hba889e8b),
	.w5(32'hbb8b5f50),
	.w6(32'h3b1f6d4b),
	.w7(32'hbaf92bd3),
	.w8(32'hbb5d3297),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a816d2f),
	.w1(32'h3b968127),
	.w2(32'hbb2ebaf9),
	.w3(32'hb9cda80d),
	.w4(32'h3c170e0d),
	.w5(32'hbad41257),
	.w6(32'h3b94e1a7),
	.w7(32'h3af96fb0),
	.w8(32'hbb273a34),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe982d3),
	.w1(32'hbab01acb),
	.w2(32'h3b31cdb1),
	.w3(32'hbb58874a),
	.w4(32'hba91980a),
	.w5(32'h3aea4ee3),
	.w6(32'h3b016c83),
	.w7(32'h3aa9ecfe),
	.w8(32'hbae7a2ce),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbace0de1),
	.w1(32'h3b64cd0f),
	.w2(32'h3930e61a),
	.w3(32'hbb02d3eb),
	.w4(32'h3b473bfb),
	.w5(32'hbbd8cf79),
	.w6(32'hba3a85f9),
	.w7(32'hbacf087d),
	.w8(32'hbb882872),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf0b645),
	.w1(32'h3ba35704),
	.w2(32'h3a9043da),
	.w3(32'hbb8826a9),
	.w4(32'h3bc1b605),
	.w5(32'h3b0e834f),
	.w6(32'h3ab41bb7),
	.w7(32'hb9e0276c),
	.w8(32'h3b8dd5a9),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4590fd),
	.w1(32'h3bddbd68),
	.w2(32'h3bcdb078),
	.w3(32'h3b938bbd),
	.w4(32'h3bcd326d),
	.w5(32'hb97b5ff0),
	.w6(32'h3b487dd3),
	.w7(32'h3bd7e01d),
	.w8(32'h39e2ae2c),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbe6bcc),
	.w1(32'h3c4c427a),
	.w2(32'hbc1ed55d),
	.w3(32'h3b10f535),
	.w4(32'hba4bef43),
	.w5(32'h3a7196c5),
	.w6(32'h3ca30bca),
	.w7(32'hbba56abd),
	.w8(32'hba2fc835),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bb226c),
	.w1(32'hbaccca8f),
	.w2(32'h3ab5ea6d),
	.w3(32'h3b304106),
	.w4(32'h3b7e9a9a),
	.w5(32'hbb995907),
	.w6(32'h3b8e5b4d),
	.w7(32'h3c4d1c8f),
	.w8(32'hba8fad5b),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeae157),
	.w1(32'hbb473139),
	.w2(32'h3ac2fd30),
	.w3(32'hbabbecdd),
	.w4(32'hbab2820d),
	.w5(32'h3a2c6252),
	.w6(32'h3abc5661),
	.w7(32'hb9aa1d37),
	.w8(32'hba596e11),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39947e94),
	.w1(32'hbb25a617),
	.w2(32'hbb3f3413),
	.w3(32'h3a2ca231),
	.w4(32'h39afeae4),
	.w5(32'h3974d65a),
	.w6(32'h3b139b82),
	.w7(32'h3aacb7e8),
	.w8(32'hb983b094),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39599f75),
	.w1(32'h3b6c43da),
	.w2(32'h3a92c0e5),
	.w3(32'h3b7844b5),
	.w4(32'h3be25c2c),
	.w5(32'h3b7f4c73),
	.w6(32'h3b42975c),
	.w7(32'hbac073db),
	.w8(32'hbaa2f883),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ba347f),
	.w1(32'h3c4e0570),
	.w2(32'h3b9f54a4),
	.w3(32'h3a80d582),
	.w4(32'h3b7eb3fa),
	.w5(32'hbb8335dc),
	.w6(32'h3c17bac9),
	.w7(32'h3c73b190),
	.w8(32'h3b8cb4fe),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b278424),
	.w1(32'hbbe63675),
	.w2(32'hbc2e0d00),
	.w3(32'h3ad10e0e),
	.w4(32'hbbbf77a7),
	.w5(32'hb9c12702),
	.w6(32'h3b659429),
	.w7(32'hbb51fe44),
	.w8(32'h3928d5e4),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a376067),
	.w1(32'hbb01909a),
	.w2(32'h39ad9ccf),
	.w3(32'h3b3f99ee),
	.w4(32'h3be52d94),
	.w5(32'hbc48bda9),
	.w6(32'hbb2b31a1),
	.w7(32'h3ba41167),
	.w8(32'hbc134e43),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4a787c),
	.w1(32'hbc913a35),
	.w2(32'hbab90078),
	.w3(32'hbba16765),
	.w4(32'hbc72a6fd),
	.w5(32'hbc11c344),
	.w6(32'hbc283005),
	.w7(32'h3a8625fa),
	.w8(32'h3b638cf3),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1306d1),
	.w1(32'hbb2036cd),
	.w2(32'hb7b30181),
	.w3(32'h3bd16dbe),
	.w4(32'hba69d299),
	.w5(32'hba52d358),
	.w6(32'hbaf335f6),
	.w7(32'hba049614),
	.w8(32'hbb07d01d),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa6f49a),
	.w1(32'h3bf9df7a),
	.w2(32'h3b9aed02),
	.w3(32'hbaf27767),
	.w4(32'h3bc48b8b),
	.w5(32'h3c07b703),
	.w6(32'h3bad7675),
	.w7(32'hb9dbd521),
	.w8(32'h3abd2a0e),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b99bcd9),
	.w1(32'hbc85c3d5),
	.w2(32'hbcac5c59),
	.w3(32'h3b4bee56),
	.w4(32'hbbce8295),
	.w5(32'hbca558e8),
	.w6(32'hbc47db7e),
	.w7(32'hb70467b5),
	.w8(32'h3b258843),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393e19b2),
	.w1(32'h3bbf474d),
	.w2(32'hbc3749e0),
	.w3(32'hbc19e1e9),
	.w4(32'hb906683f),
	.w5(32'h3b4863a1),
	.w6(32'h3b9b75ba),
	.w7(32'hbbb3545b),
	.w8(32'hbb3db85b),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1018bf),
	.w1(32'h3ac86311),
	.w2(32'hba6a152f),
	.w3(32'hbba11819),
	.w4(32'h3a8b1d54),
	.w5(32'h3a9788a9),
	.w6(32'h39d03d11),
	.w7(32'hba18bc6c),
	.w8(32'h3928822f),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aae43b1),
	.w1(32'h3b1b00ab),
	.w2(32'hbb68cfbd),
	.w3(32'h3a65897d),
	.w4(32'h3bc0612a),
	.w5(32'h39d78e9b),
	.w6(32'h3b3847d4),
	.w7(32'h3b225543),
	.w8(32'h3b08528d),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule