module layer_10_featuremap_281(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb53c351b),
	.w1(32'hb68aa357),
	.w2(32'hb6bfec84),
	.w3(32'hb7935a06),
	.w4(32'hb712eac3),
	.w5(32'h35a15188),
	.w6(32'hb78ca76a),
	.w7(32'hb71626ec),
	.w8(32'h370151ec),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36d580e6),
	.w1(32'hb712f7e0),
	.w2(32'hb7750bbe),
	.w3(32'hb6e501d1),
	.w4(32'hb6b01e7d),
	.w5(32'h36a77372),
	.w6(32'hb5e343f6),
	.w7(32'h36e84197),
	.w8(32'hb6afc6ad),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb74c36d7),
	.w1(32'hb8346d4a),
	.w2(32'hb7b77b40),
	.w3(32'hb826e86d),
	.w4(32'hb773eac5),
	.w5(32'hb617d60f),
	.w6(32'hb83a5227),
	.w7(32'hb7927d6a),
	.w8(32'hb3e2414b),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h360af29c),
	.w1(32'h370dcb7d),
	.w2(32'hb60545ac),
	.w3(32'h3605d1ef),
	.w4(32'hb7233460),
	.w5(32'h37beb689),
	.w6(32'h375ed86d),
	.w7(32'h35b1427d),
	.w8(32'h35ed6c2e),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38117a07),
	.w1(32'h380dd9d3),
	.w2(32'hb5db7db1),
	.w3(32'h383a38f5),
	.w4(32'h37b8c779),
	.w5(32'hb6c0a5a1),
	.w6(32'h379037d8),
	.w7(32'hb7347261),
	.w8(32'hb684479b),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35f3d47e),
	.w1(32'h36256311),
	.w2(32'hb68c072d),
	.w3(32'h345fa311),
	.w4(32'h36697b21),
	.w5(32'h35a14998),
	.w6(32'h35d9a366),
	.w7(32'h3386bfd1),
	.w8(32'hb3959c21),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb4044ff1),
	.w1(32'hb556a1e4),
	.w2(32'hb6da6671),
	.w3(32'h37135867),
	.w4(32'hb69b1514),
	.w5(32'h37747efc),
	.w6(32'h3738ad65),
	.w7(32'hb67aa66e),
	.w8(32'h36bc146b),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h366d37dd),
	.w1(32'h382e5b3d),
	.w2(32'h37e16efc),
	.w3(32'h38012f21),
	.w4(32'h36eb87b1),
	.w5(32'h370ed67c),
	.w6(32'h36efbec8),
	.w7(32'h37cfbbf4),
	.w8(32'h359233b9),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7643a0d),
	.w1(32'h3779180c),
	.w2(32'h37e8106b),
	.w3(32'hb8055cdc),
	.w4(32'h36e123b1),
	.w5(32'h373ce38f),
	.w6(32'hb84ee0a9),
	.w7(32'hb7fe4f32),
	.w8(32'h36aa60ce),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38126c07),
	.w1(32'h3893a5b9),
	.w2(32'h393060a2),
	.w3(32'hb8cf1ae1),
	.w4(32'hb81c3a8d),
	.w5(32'h39046c82),
	.w6(32'hb8938ab9),
	.w7(32'hb8942870),
	.w8(32'h35348924),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb86a2b70),
	.w1(32'hb7f60a36),
	.w2(32'hb85a1cbe),
	.w3(32'hb7904fc3),
	.w4(32'h3749c9ce),
	.w5(32'h36cbedd1),
	.w6(32'hb8199110),
	.w7(32'h36d4984a),
	.w8(32'h376cd547),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb765915d),
	.w1(32'hb76d07f5),
	.w2(32'hb85fb674),
	.w3(32'h3740f0d5),
	.w4(32'hb65a85e3),
	.w5(32'hb7d52109),
	.w6(32'h3796b19b),
	.w7(32'h3800f354),
	.w8(32'hb7303fe3),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h374eb0b4),
	.w1(32'h36aa2b68),
	.w2(32'h3860caa1),
	.w3(32'hb7fefae4),
	.w4(32'hb8608ec9),
	.w5(32'h3837bf50),
	.w6(32'hb835c299),
	.w7(32'hb8987abe),
	.w8(32'hb74524ed),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8797185),
	.w1(32'hb87bf23a),
	.w2(32'hb88c01b7),
	.w3(32'h378afa5e),
	.w4(32'hb769de5c),
	.w5(32'hb821491b),
	.w6(32'h38518765),
	.w7(32'hb71eb5c9),
	.w8(32'hb7d2dc2e),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb75f42cf),
	.w1(32'h3858aef3),
	.w2(32'h390b3034),
	.w3(32'hb93aa123),
	.w4(32'hb8e52acc),
	.w5(32'hb7429abc),
	.w6(32'hb8af9388),
	.w7(32'hb8fd31b7),
	.w8(32'hb8a7660b),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7f3ce2d),
	.w1(32'h38b04652),
	.w2(32'h3918785e),
	.w3(32'hb8925d4b),
	.w4(32'h384b5a79),
	.w5(32'h38c3b87a),
	.w6(32'hb81d66f9),
	.w7(32'hb72de506),
	.w8(32'h37dff4b2),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36d1e6e7),
	.w1(32'h37779f77),
	.w2(32'hb64956d6),
	.w3(32'h359433ad),
	.w4(32'h384e705f),
	.w5(32'h381b68c9),
	.w6(32'hb81a536d),
	.w7(32'h37a1346d),
	.w8(32'h37d292c8),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35e560d4),
	.w1(32'hb705591b),
	.w2(32'h3887dcf9),
	.w3(32'hb7301cdd),
	.w4(32'hb6316185),
	.w5(32'h388dccd4),
	.w6(32'hb818f86e),
	.w7(32'hb883c300),
	.w8(32'hb7181d26),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h371ce9ee),
	.w1(32'h37b8054d),
	.w2(32'h37ac69c4),
	.w3(32'h363186eb),
	.w4(32'h38506fe7),
	.w5(32'h38849767),
	.w6(32'hb8117c3d),
	.w7(32'hb7d9fba4),
	.w8(32'h37b01b43),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7812968),
	.w1(32'hb7c4d093),
	.w2(32'hb7526a32),
	.w3(32'h3708ac18),
	.w4(32'hb5b59c0a),
	.w5(32'hb3fc53a2),
	.w6(32'hb7903588),
	.w7(32'hb776127c),
	.w8(32'hb6bef635),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6218104),
	.w1(32'h37d37735),
	.w2(32'h38143acd),
	.w3(32'h380f1b77),
	.w4(32'h37e94197),
	.w5(32'hb7693708),
	.w6(32'h38496d13),
	.w7(32'h383aad1f),
	.w8(32'hb6e63dd1),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7b60330),
	.w1(32'h3742a351),
	.w2(32'hb7a499fc),
	.w3(32'hb6799ef8),
	.w4(32'h373d1db5),
	.w5(32'hb67db1b7),
	.w6(32'h37a5396c),
	.w7(32'h37f30628),
	.w8(32'h3730be8d),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389409b3),
	.w1(32'hb8155563),
	.w2(32'h39005c8f),
	.w3(32'hb84c231c),
	.w4(32'hb9252936),
	.w5(32'h376aaf68),
	.w6(32'hb85c49d0),
	.w7(32'hb91b79cd),
	.w8(32'hb88b7109),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35abe578),
	.w1(32'h389c2092),
	.w2(32'h38d4a8cb),
	.w3(32'hb8009c78),
	.w4(32'hb7965810),
	.w5(32'h384deaf9),
	.w6(32'h37b508d7),
	.w7(32'hb8750e1e),
	.w8(32'hb79d01fe),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb4b12a88),
	.w1(32'h3761da6d),
	.w2(32'h3758e880),
	.w3(32'hb6d92207),
	.w4(32'h36c68253),
	.w5(32'hb73e1bca),
	.w6(32'hb885cae7),
	.w7(32'hb75cc72e),
	.w8(32'hb7002f2e),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3507c155),
	.w1(32'hb791ad72),
	.w2(32'h37c4a057),
	.w3(32'hb860b173),
	.w4(32'hb84b3767),
	.w5(32'h3793c3b5),
	.w6(32'hb8178b05),
	.w7(32'hb7da6f03),
	.w8(32'hb7840223),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h34bb2229),
	.w1(32'hb7013f36),
	.w2(32'hb69014cf),
	.w3(32'hb558b9b4),
	.w4(32'hb7683d1f),
	.w5(32'hb782a469),
	.w6(32'hb77c79f5),
	.w7(32'hb701d168),
	.w8(32'hb79b6df2),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7daa02b),
	.w1(32'hb791d77e),
	.w2(32'hb7e3e2aa),
	.w3(32'hb75c7f59),
	.w4(32'h3786394d),
	.w5(32'hb775ab5b),
	.w6(32'hb7f5e6f4),
	.w7(32'hb64e9604),
	.w8(32'hb7261a79),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7c4a062),
	.w1(32'h35ec7cf7),
	.w2(32'hb735f042),
	.w3(32'hb7322a2c),
	.w4(32'h3758b6ff),
	.w5(32'h37848f9b),
	.w6(32'hb7574cf9),
	.w7(32'h381440ca),
	.w8(32'h3822df38),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36f84f1f),
	.w1(32'h37d6aaad),
	.w2(32'h38f473b5),
	.w3(32'hb8be049e),
	.w4(32'hb87861fd),
	.w5(32'h388e414b),
	.w6(32'hb857ea45),
	.w7(32'hb8a30535),
	.w8(32'hb7ce5144),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb60bfdac),
	.w1(32'hb7ab367d),
	.w2(32'hb6e1bf87),
	.w3(32'h3703fb19),
	.w4(32'hb72c4f57),
	.w5(32'h378dc644),
	.w6(32'hb82652ae),
	.w7(32'hb834e816),
	.w8(32'hb5caa710),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb82d139b),
	.w1(32'h36147384),
	.w2(32'hb7718822),
	.w3(32'hb79e7a98),
	.w4(32'hb69b27bc),
	.w5(32'h37181286),
	.w6(32'hb7958be9),
	.w7(32'h3654bc6f),
	.w8(32'h37939dfc),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h369aae74),
	.w1(32'h3808ae88),
	.w2(32'h38a14029),
	.w3(32'hb7d3f62b),
	.w4(32'hb75aaf11),
	.w5(32'h3848cbc5),
	.w6(32'hb814e837),
	.w7(32'hb88c2822),
	.w8(32'hb64e916e),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37d45654),
	.w1(32'h37dc4bde),
	.w2(32'h3846e0d9),
	.w3(32'h378f66b7),
	.w4(32'h380c4375),
	.w5(32'h385f014a),
	.w6(32'hb7ec0023),
	.w7(32'hb79da320),
	.w8(32'h374f85a5),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3701c09b),
	.w1(32'h374e9bcd),
	.w2(32'h379d55cb),
	.w3(32'h36773fff),
	.w4(32'h36af836e),
	.w5(32'hb565feae),
	.w6(32'hb79f3a34),
	.w7(32'h3654ba2b),
	.w8(32'hb74a2001),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb4f6bf50),
	.w1(32'hb4fc63db),
	.w2(32'hb71dc0af),
	.w3(32'h36885506),
	.w4(32'hb7384e77),
	.w5(32'hb7451ca0),
	.w6(32'h36112d60),
	.w7(32'hb7f475d4),
	.w8(32'h35e2208a),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h372775e2),
	.w1(32'hb90dd54b),
	.w2(32'hb7e92079),
	.w3(32'hb7981edc),
	.w4(32'hb928f6d8),
	.w5(32'hb6803a67),
	.w6(32'hb8565765),
	.w7(32'hb9122cba),
	.w8(32'hb80fb9ac),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8117849),
	.w1(32'hb76c0081),
	.w2(32'hb881b287),
	.w3(32'h38a985f4),
	.w4(32'h386f9df2),
	.w5(32'hb8272b86),
	.w6(32'h389908f9),
	.w7(32'h387ffe2f),
	.w8(32'h37f5f5cc),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb810aefe),
	.w1(32'hb666fcdd),
	.w2(32'hb8f4b87b),
	.w3(32'h37aa8b13),
	.w4(32'h3884606b),
	.w5(32'hb8442598),
	.w6(32'h36a0f8cd),
	.w7(32'h38846724),
	.w8(32'h37cfce2b),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h381849ae),
	.w1(32'h384f1e96),
	.w2(32'h37c4dc51),
	.w3(32'h383f4ff8),
	.w4(32'h38287d20),
	.w5(32'h379a8dd9),
	.w6(32'h3873cd34),
	.w7(32'h3817e221),
	.w8(32'h37bc220d),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37c39c46),
	.w1(32'h3675a8a3),
	.w2(32'h36e4ed67),
	.w3(32'h37429172),
	.w4(32'h37d08165),
	.w5(32'h3591feef),
	.w6(32'h378947eb),
	.w7(32'h37ad79a9),
	.w8(32'h3609fc00),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36daf6ab),
	.w1(32'h3717c376),
	.w2(32'h35b4d209),
	.w3(32'h3344a644),
	.w4(32'hb6a4607d),
	.w5(32'h377e9bd3),
	.w6(32'h36321335),
	.w7(32'h3692cf05),
	.w8(32'hb6dc309b),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37564561),
	.w1(32'h363298aa),
	.w2(32'hb712db52),
	.w3(32'h37b42c5f),
	.w4(32'h37127789),
	.w5(32'h37e6fdba),
	.w6(32'hb71ae925),
	.w7(32'hb806f90d),
	.w8(32'h36bc4dc4),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a9c6c2),
	.w1(32'h3801a7e8),
	.w2(32'h3920fa93),
	.w3(32'hb9227131),
	.w4(32'hb6dcd33d),
	.w5(32'h38c66c0f),
	.w6(32'hb91c7818),
	.w7(32'hb8d1ee83),
	.w8(32'hb7bf2a3d),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6cd7767),
	.w1(32'h383b6502),
	.w2(32'h390f552b),
	.w3(32'hb81479b4),
	.w4(32'hb7175814),
	.w5(32'h3894b663),
	.w6(32'hb889a2b4),
	.w7(32'hb88f5a4c),
	.w8(32'hb745e535),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36bd94d0),
	.w1(32'h38162706),
	.w2(32'h39149924),
	.w3(32'hb8a7eb95),
	.w4(32'hb80a4d8c),
	.w5(32'h389900de),
	.w6(32'hb8d0c577),
	.w7(32'hb892d5c7),
	.w8(32'hb716b85d),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h378d79e9),
	.w1(32'h3843c4af),
	.w2(32'h38f95b78),
	.w3(32'h33990e61),
	.w4(32'h37d4d6d8),
	.w5(32'h38616648),
	.w6(32'hb7ab4c8a),
	.w7(32'hb7427859),
	.w8(32'hb6a8e91d),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3457ed82),
	.w1(32'h37bcecb8),
	.w2(32'hb7947d32),
	.w3(32'hb8115b93),
	.w4(32'hb85664cb),
	.w5(32'h37a6cb05),
	.w6(32'hb811a90b),
	.w7(32'hb81a636c),
	.w8(32'hb7691d75),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6d45563),
	.w1(32'h3732ddf1),
	.w2(32'h378cebbd),
	.w3(32'h3426bac8),
	.w4(32'h3727697c),
	.w5(32'hb70dc82d),
	.w6(32'h34d0f46d),
	.w7(32'hb5e1160d),
	.w8(32'hb773551d),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36ab8896),
	.w1(32'h38d951c9),
	.w2(32'h38bb4e0a),
	.w3(32'hb7bd5227),
	.w4(32'h388228d0),
	.w5(32'h38c0aec2),
	.w6(32'hb858e920),
	.w7(32'hb78099e7),
	.w8(32'h3810058f),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h372a6fbe),
	.w1(32'hb5f7856d),
	.w2(32'hb4c1bdb7),
	.w3(32'h362d0134),
	.w4(32'hb557362c),
	.w5(32'h38286110),
	.w6(32'h371ee760),
	.w7(32'hb7b653ae),
	.w8(32'h378822cb),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h378f2c1c),
	.w1(32'h3747e7ce),
	.w2(32'h378c8d75),
	.w3(32'h37d34132),
	.w4(32'h3703c67f),
	.w5(32'h36248b27),
	.w6(32'h379f2388),
	.w7(32'h352dee4d),
	.w8(32'h366293b6),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37b3303b),
	.w1(32'h37e9cc76),
	.w2(32'h369445ea),
	.w3(32'h3780fbd2),
	.w4(32'h37daab7c),
	.w5(32'h37b2f738),
	.w6(32'hb7929c86),
	.w7(32'hb7bd69dc),
	.w8(32'h37a13f2a),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38aac4b0),
	.w1(32'h38bc9fc6),
	.w2(32'h38e036a7),
	.w3(32'hb729f0fd),
	.w4(32'h3627681c),
	.w5(32'h39267a2d),
	.w6(32'hb8c9316e),
	.w7(32'hb8e7eff8),
	.w8(32'h37b6a2f9),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h372aa55a),
	.w1(32'h378964bf),
	.w2(32'h373f8851),
	.w3(32'h37b81292),
	.w4(32'h37bfa80d),
	.w5(32'h370dea2d),
	.w6(32'h367e2512),
	.w7(32'h36923458),
	.w8(32'hb74534ac),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6e9704f),
	.w1(32'hb49b388f),
	.w2(32'h37345bf0),
	.w3(32'h37d44681),
	.w4(32'h37bb4d28),
	.w5(32'h362f257a),
	.w6(32'hb5516af4),
	.w7(32'h36cac47a),
	.w8(32'hb5fb4afa),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h364798e0),
	.w1(32'hb726be29),
	.w2(32'h3683ea60),
	.w3(32'h36e65733),
	.w4(32'h3789b033),
	.w5(32'hb685f7eb),
	.w6(32'hb608418d),
	.w7(32'h35eb2de6),
	.w8(32'hb76dc4b4),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb427e50a),
	.w1(32'hb8132f84),
	.w2(32'hb7af6540),
	.w3(32'hb80f0d84),
	.w4(32'hb76e6e89),
	.w5(32'hb736fd20),
	.w6(32'hb801cdc9),
	.w7(32'hb7a31aeb),
	.w8(32'hb6ffbaa9),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6f882d2),
	.w1(32'h37e5d6f2),
	.w2(32'hb75d7eef),
	.w3(32'h36fabdc5),
	.w4(32'h3632e9b1),
	.w5(32'h36ab1762),
	.w6(32'h372c07f0),
	.w7(32'h362436fa),
	.w8(32'hb7458ffa),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb782b86f),
	.w1(32'hb6fd3822),
	.w2(32'hb6b40dc1),
	.w3(32'hb4f5d134),
	.w4(32'h37a97e06),
	.w5(32'hb7a82ffd),
	.w6(32'hb870a754),
	.w7(32'hb7e41911),
	.w8(32'h36358cd6),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb70be184),
	.w1(32'h381f81e5),
	.w2(32'h382bef6f),
	.w3(32'hb898378e),
	.w4(32'h3809bc6a),
	.w5(32'h382e399b),
	.w6(32'hb8809f54),
	.w7(32'hb7ae6869),
	.w8(32'h37a9702e),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37cca8d4),
	.w1(32'h373cfd6b),
	.w2(32'h37caff61),
	.w3(32'hb58ab5d5),
	.w4(32'h36178513),
	.w5(32'h3411e561),
	.w6(32'hb6350617),
	.w7(32'h373c70a1),
	.w8(32'hb7ff9844),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37756b0a),
	.w1(32'h37299ac3),
	.w2(32'h37acf932),
	.w3(32'h3763c0a7),
	.w4(32'h3795b2fc),
	.w5(32'h3751e234),
	.w6(32'hb81ac23b),
	.w7(32'hb7990a67),
	.w8(32'h3727d225),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h371d609e),
	.w1(32'h36529162),
	.w2(32'h373d76f9),
	.w3(32'h3768ce93),
	.w4(32'h37788e68),
	.w5(32'h372460c1),
	.w6(32'h37169d6c),
	.w7(32'h3726efdf),
	.w8(32'h3712dc34),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36fca817),
	.w1(32'h356752b5),
	.w2(32'h3759197d),
	.w3(32'hb6866570),
	.w4(32'h37296109),
	.w5(32'h3746c472),
	.w6(32'h36b549bb),
	.w7(32'h3699793a),
	.w8(32'hb6b7363b),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3789ad60),
	.w1(32'h371dd021),
	.w2(32'h36a641aa),
	.w3(32'h3748fcea),
	.w4(32'h37e00e81),
	.w5(32'h36bda41a),
	.w6(32'hb7fcc8a5),
	.w7(32'hb6e83676),
	.w8(32'h36eb9bfa),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3730d816),
	.w1(32'h37553f26),
	.w2(32'hb62acea5),
	.w3(32'hb727b705),
	.w4(32'hb79a98df),
	.w5(32'h38395f9c),
	.w6(32'hb700eeae),
	.w7(32'hb7b15794),
	.w8(32'h37b741b9),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h374e0409),
	.w1(32'h35fa1086),
	.w2(32'h37418636),
	.w3(32'hb82ab1a5),
	.w4(32'hb812ca29),
	.w5(32'h37f101a3),
	.w6(32'hb82694a2),
	.w7(32'hb866cf63),
	.w8(32'h358c6e8a),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb693c39b),
	.w1(32'h36d9e1ad),
	.w2(32'hb78b9354),
	.w3(32'hb6355b2e),
	.w4(32'h3721baca),
	.w5(32'h37010c55),
	.w6(32'h3765efc5),
	.w7(32'h374ed460),
	.w8(32'h378399aa),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb75adbaa),
	.w1(32'hb804c3f5),
	.w2(32'h36af7404),
	.w3(32'hb85846db),
	.w4(32'hb8bae2b5),
	.w5(32'hb761bf3e),
	.w6(32'hb80fd699),
	.w7(32'hb8bf9f12),
	.w8(32'hb84e1797),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36b3848f),
	.w1(32'hb76b20f3),
	.w2(32'hb6a6bc06),
	.w3(32'h36cecb0a),
	.w4(32'hb6a8a1a1),
	.w5(32'hb7ac7244),
	.w6(32'hb804bb9b),
	.w7(32'hb7e73ca9),
	.w8(32'hb74fb96a),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37414270),
	.w1(32'h380051a7),
	.w2(32'h378b88c3),
	.w3(32'hb7587643),
	.w4(32'h37b14e29),
	.w5(32'hb7148388),
	.w6(32'h37de71e7),
	.w7(32'h3842bdee),
	.w8(32'h37326f91),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37ee014e),
	.w1(32'h37349a24),
	.w2(32'hb73da8b4),
	.w3(32'hb7aabf9d),
	.w4(32'hb71d974f),
	.w5(32'h3753e40f),
	.w6(32'hb68ecd61),
	.w7(32'h36f3a217),
	.w8(32'h37343665),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3592d988),
	.w1(32'hb748e979),
	.w2(32'hb7b20e13),
	.w3(32'h37115ae0),
	.w4(32'h365d7ced),
	.w5(32'h3544a5ae),
	.w6(32'hb786540e),
	.w7(32'h36814486),
	.w8(32'h36bd98b3),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h342287e2),
	.w1(32'hb603aede),
	.w2(32'hb7b82149),
	.w3(32'h34c6c901),
	.w4(32'hb78e4738),
	.w5(32'h379abd5d),
	.w6(32'h36dbe0b8),
	.w7(32'hb7ccaa31),
	.w8(32'h371288a8),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37401caa),
	.w1(32'h36e79012),
	.w2(32'h37514799),
	.w3(32'h374b496d),
	.w4(32'h3757f9fc),
	.w5(32'h374cb2b0),
	.w6(32'h374af039),
	.w7(32'h36ec256b),
	.w8(32'hb70f4b45),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a3c84c),
	.w1(32'h3837673c),
	.w2(32'h38c8606c),
	.w3(32'hb8d8adc6),
	.w4(32'h385813be),
	.w5(32'h37e13ddb),
	.w6(32'hb86517e3),
	.w7(32'h37692871),
	.w8(32'h369fec85),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7ec886f),
	.w1(32'hb7546133),
	.w2(32'h3781cb49),
	.w3(32'hb7ab7b8f),
	.w4(32'h353c7f9b),
	.w5(32'hb6f62343),
	.w6(32'hb7db71e6),
	.w7(32'hb7e7fd5b),
	.w8(32'hb76f3636),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7dbe944),
	.w1(32'hb84e1fa6),
	.w2(32'hb882b9e4),
	.w3(32'hb7fbde6a),
	.w4(32'hb88b3d28),
	.w5(32'hb8445bbc),
	.w6(32'h36f84576),
	.w7(32'hb82f032c),
	.w8(32'hb828c862),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36fb13d3),
	.w1(32'hb685e847),
	.w2(32'hb66f8997),
	.w3(32'hb7c45e35),
	.w4(32'hb755bf96),
	.w5(32'hb779d9dd),
	.w6(32'hb7aba8db),
	.w7(32'hb7112834),
	.w8(32'h353d3772),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb791f789),
	.w1(32'h35e445ee),
	.w2(32'h385c8803),
	.w3(32'hb89453bf),
	.w4(32'hb8945adb),
	.w5(32'h38245926),
	.w6(32'hb7caffda),
	.w7(32'hb87f1e2d),
	.w8(32'hb7b23dd2),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37727230),
	.w1(32'hb72df465),
	.w2(32'hb784a1e5),
	.w3(32'h373f478b),
	.w4(32'h37c2a46d),
	.w5(32'hb6f1901d),
	.w6(32'hb730583b),
	.w7(32'hb6f03d1a),
	.w8(32'hb6d75b06),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb65c7dcb),
	.w1(32'hb7cf4d57),
	.w2(32'hb7199046),
	.w3(32'hb8011500),
	.w4(32'hb797913e),
	.w5(32'hb80641ec),
	.w6(32'hb6d00620),
	.w7(32'hb6e0c52d),
	.w8(32'hb7e78a3f),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6a7fab9),
	.w1(32'h36b1a3c0),
	.w2(32'hb7921970),
	.w3(32'hb7ee3286),
	.w4(32'hb8395daa),
	.w5(32'h36db490a),
	.w6(32'h37345267),
	.w7(32'hb7fc8bb5),
	.w8(32'hb73488bd),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb745f767),
	.w1(32'hb7d289df),
	.w2(32'hb75bc776),
	.w3(32'hb6e590c6),
	.w4(32'hb63c0efd),
	.w5(32'h364dd5c8),
	.w6(32'hb7687ab3),
	.w7(32'hb572458b),
	.w8(32'hb69e7e58),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb735c559),
	.w1(32'hb7d5dd79),
	.w2(32'h3793824e),
	.w3(32'hb7987815),
	.w4(32'h36bfea56),
	.w5(32'h36bf2251),
	.w6(32'hb824e398),
	.w7(32'h3734bfb7),
	.w8(32'h360f20ee),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37755636),
	.w1(32'hb81424a0),
	.w2(32'hb813ca66),
	.w3(32'hb7becf4b),
	.w4(32'hb7d454c1),
	.w5(32'h377c27cc),
	.w6(32'hb7fcbb41),
	.w7(32'hb748dd0d),
	.w8(32'hb6d54b91),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6da9991),
	.w1(32'hb75f3625),
	.w2(32'hb7883b3c),
	.w3(32'h377e59c6),
	.w4(32'h37bcd36b),
	.w5(32'hb6fd4c04),
	.w6(32'hb81c83f0),
	.w7(32'hb6e55c11),
	.w8(32'hb65352fd),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h381ecd6d),
	.w1(32'h374a8aa7),
	.w2(32'h3823ba90),
	.w3(32'hb625fd17),
	.w4(32'hb73d4a7a),
	.w5(32'h3862a878),
	.w6(32'hb7e67016),
	.w7(32'hb7eb9624),
	.w8(32'h371a109e),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6b55b65),
	.w1(32'h36e8bc25),
	.w2(32'h37b3b2c4),
	.w3(32'hb7aa78d2),
	.w4(32'h37aef661),
	.w5(32'hb7094209),
	.w6(32'h37b80a1c),
	.w7(32'h382e5908),
	.w8(32'h3751adc9),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb78bcc02),
	.w1(32'h37c53fa5),
	.w2(32'hb8773aa5),
	.w3(32'h3813476c),
	.w4(32'hb7897d52),
	.w5(32'hb83e63c2),
	.w6(32'h3896f886),
	.w7(32'hb69c5a0d),
	.w8(32'hb81b4f8f),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37de8682),
	.w1(32'h380b42a0),
	.w2(32'h3907476e),
	.w3(32'hb8b7c24b),
	.w4(32'hb6c31279),
	.w5(32'h390def9c),
	.w6(32'hb8c0d142),
	.w7(32'hb8b57eeb),
	.w8(32'hb85eeda9),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8318534),
	.w1(32'hb7a4ef3f),
	.w2(32'hb89196ef),
	.w3(32'h382182c9),
	.w4(32'h3784e790),
	.w5(32'hb7c44c80),
	.w6(32'h353a6fd0),
	.w7(32'h369a16e2),
	.w8(32'hb7a6189d),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb79eeec7),
	.w1(32'hb810ca61),
	.w2(32'h38ca18b0),
	.w3(32'hb9306589),
	.w4(32'hb8231620),
	.w5(32'h37b9f918),
	.w6(32'hb938aec2),
	.w7(32'hb8adde24),
	.w8(32'hb7c70b4f),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb68490fd),
	.w1(32'h38a5d4b0),
	.w2(32'h39036eb1),
	.w3(32'hb8c4f9c3),
	.w4(32'hb7dc5641),
	.w5(32'h3901a852),
	.w6(32'hb8e73d68),
	.w7(32'hb8a75deb),
	.w8(32'h36978809),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6f5f088),
	.w1(32'h37b35dbc),
	.w2(32'h37ea483c),
	.w3(32'hb79caa74),
	.w4(32'hb6d70f65),
	.w5(32'hb771bdf9),
	.w6(32'hb7c68efc),
	.w7(32'hb7b7a000),
	.w8(32'hb79997b2),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb83765e9),
	.w1(32'hb7e73093),
	.w2(32'hb8383ee2),
	.w3(32'h34f89eea),
	.w4(32'h35f318c7),
	.w5(32'hb6bacf6a),
	.w6(32'hb7984383),
	.w7(32'hb7949c3c),
	.w8(32'hb73b5108),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3710fc9a),
	.w1(32'h3882465a),
	.w2(32'h39357a58),
	.w3(32'hb8879036),
	.w4(32'hb7bf4eec),
	.w5(32'h3bbf5548),
	.w6(32'hb8a9a3a1),
	.w7(32'hb90eb66c),
	.w8(32'h3c07b837),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf12ce3),
	.w1(32'h3bcbdb10),
	.w2(32'h3bb8c61b),
	.w3(32'h3b79b2c6),
	.w4(32'h3b1e3e29),
	.w5(32'hba980145),
	.w6(32'h3c1caff9),
	.w7(32'h3bbe5988),
	.w8(32'hbbb7262c),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe98b3c),
	.w1(32'hbba9ea7e),
	.w2(32'hbbe6500d),
	.w3(32'hbba53193),
	.w4(32'hbb55b8bd),
	.w5(32'hbb9d258b),
	.w6(32'hbb6c5007),
	.w7(32'hbb511d88),
	.w8(32'h3ba415b0),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaecef6d),
	.w1(32'h3b407c67),
	.w2(32'hbb55dcae),
	.w3(32'hbba66746),
	.w4(32'hbc0aaaad),
	.w5(32'h3bbd8dd3),
	.w6(32'h3c9fe94b),
	.w7(32'h3be9cac8),
	.w8(32'hbb1096cc),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c544d86),
	.w1(32'h3ca4c4eb),
	.w2(32'h3cae4bf8),
	.w3(32'h3bd3f46c),
	.w4(32'h3baeeb66),
	.w5(32'hbb65c4c6),
	.w6(32'hbb4ebf5a),
	.w7(32'h3a5015e0),
	.w8(32'hbc19128d),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9df13a),
	.w1(32'h3b70f981),
	.w2(32'h3b57ac25),
	.w3(32'hbbde9b49),
	.w4(32'hbb42d4ec),
	.w5(32'h3b315c3e),
	.w6(32'hbbb23acd),
	.w7(32'h3b18d25d),
	.w8(32'h3a54459b),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb87371d),
	.w1(32'hbb4e028b),
	.w2(32'hbb86af02),
	.w3(32'hb9b402f1),
	.w4(32'hbbac1976),
	.w5(32'hba9443bc),
	.w6(32'hbbe322d8),
	.w7(32'hbb7b6bad),
	.w8(32'h3c06696d),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb21f0c0),
	.w1(32'h3bb682c1),
	.w2(32'h39bf58be),
	.w3(32'hbb055b8d),
	.w4(32'hb96802a6),
	.w5(32'h3b0480bc),
	.w6(32'h3c6cf20e),
	.w7(32'h3b99e405),
	.w8(32'hbbb9eff8),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5f261d),
	.w1(32'hbb183b9f),
	.w2(32'h3ac918cc),
	.w3(32'hba97b4d5),
	.w4(32'h3b55fbbf),
	.w5(32'hbc035e9c),
	.w6(32'hbbdb990d),
	.w7(32'hbafcce7e),
	.w8(32'hbbcf77a6),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc14b5ff),
	.w1(32'hbc1bfd71),
	.w2(32'hbc2945da),
	.w3(32'hbba62780),
	.w4(32'hbb8e90b9),
	.w5(32'h3bd34732),
	.w6(32'hbc0ce8b5),
	.w7(32'hbc09a476),
	.w8(32'h3b9873e0),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3d0de3),
	.w1(32'h3bf3ae8a),
	.w2(32'h3b573dc4),
	.w3(32'h3c1167f6),
	.w4(32'h3ba8a1c8),
	.w5(32'h3b81570d),
	.w6(32'h3c77dc2b),
	.w7(32'h3c1bebc3),
	.w8(32'h3bf928d9),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc8b937),
	.w1(32'h3bac0da4),
	.w2(32'h3bbce97a),
	.w3(32'h3b0da32d),
	.w4(32'h3a982cf3),
	.w5(32'h3b80455f),
	.w6(32'h3c2065b7),
	.w7(32'h3bbb8a3f),
	.w8(32'h3b80e44f),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9eac72),
	.w1(32'h3b411f8b),
	.w2(32'hba91caa6),
	.w3(32'h3b2bb974),
	.w4(32'hb8b0df82),
	.w5(32'hba2c2d03),
	.w6(32'h3be86bbb),
	.w7(32'hb9ffab21),
	.w8(32'hbadcc791),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9355ce),
	.w1(32'hbbb9fd49),
	.w2(32'hbbc6d376),
	.w3(32'hba608737),
	.w4(32'hba32f825),
	.w5(32'h3aae8936),
	.w6(32'hba9a935e),
	.w7(32'hbb260099),
	.w8(32'h3ad97ff7),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba994f76),
	.w1(32'hbb69ccd9),
	.w2(32'hbbbeee2c),
	.w3(32'h3b9ededd),
	.w4(32'hbb2ec951),
	.w5(32'h3b9eb307),
	.w6(32'hbc0f1400),
	.w7(32'hbc2531c9),
	.w8(32'hb8c7eac9),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3ec4ad),
	.w1(32'h3a4c1535),
	.w2(32'h3b80242c),
	.w3(32'h3986a92c),
	.w4(32'h3b564060),
	.w5(32'h3c198c10),
	.w6(32'hbb45ff06),
	.w7(32'h3a47ba75),
	.w8(32'hbad8d6b4),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c81bf9d),
	.w1(32'h3c6d43df),
	.w2(32'h3c4c22de),
	.w3(32'h3b592fc6),
	.w4(32'h3bd24ea2),
	.w5(32'hbb01930c),
	.w6(32'hbbd60271),
	.w7(32'hbb8dd62a),
	.w8(32'hbb444d1f),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8091c2),
	.w1(32'hbb9b5a86),
	.w2(32'hba4b7a69),
	.w3(32'h3b0db0f0),
	.w4(32'h3a3b1021),
	.w5(32'hbb83fee1),
	.w6(32'h3abda006),
	.w7(32'h3b241280),
	.w8(32'h3a8a65d2),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbf329f),
	.w1(32'hbb4aefca),
	.w2(32'hb99e75b7),
	.w3(32'h3b50f9a7),
	.w4(32'hbb85be4a),
	.w5(32'hba25e888),
	.w6(32'hbbd053c2),
	.w7(32'hbb9e541c),
	.w8(32'hbb2733e2),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad1de33),
	.w1(32'h3bb93b24),
	.w2(32'h3c32ce53),
	.w3(32'h3a74334a),
	.w4(32'h3bf45601),
	.w5(32'h3b4de8c2),
	.w6(32'h3afb26e5),
	.w7(32'h3c227ab2),
	.w8(32'h3bf32b35),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c096f18),
	.w1(32'h3c21622d),
	.w2(32'hbb10619f),
	.w3(32'h3aa252d6),
	.w4(32'hbb88dca0),
	.w5(32'hbb920770),
	.w6(32'hba832e62),
	.w7(32'hbb8336d9),
	.w8(32'hb9427599),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf256a5),
	.w1(32'hbc0e99dd),
	.w2(32'hbc5a9388),
	.w3(32'hbc1722f7),
	.w4(32'hbc4dbbdd),
	.w5(32'h3bd70199),
	.w6(32'hbafe36b4),
	.w7(32'hbbcf966d),
	.w8(32'h3bdbda6b),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aabc13f),
	.w1(32'h3b4fadff),
	.w2(32'hbb910d3a),
	.w3(32'h3adf805b),
	.w4(32'hbbdd6725),
	.w5(32'hbca6687f),
	.w6(32'h3b4c5b96),
	.w7(32'hbbaf2d0b),
	.w8(32'h3b99bf49),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2222e5),
	.w1(32'h3c0cf4b2),
	.w2(32'h3c028309),
	.w3(32'h3a0b47cb),
	.w4(32'hbb42ec00),
	.w5(32'h3a4dea48),
	.w6(32'h3cb76671),
	.w7(32'h3c89f60b),
	.w8(32'h3a2f8122),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac92203),
	.w1(32'hba610e95),
	.w2(32'hbb037415),
	.w3(32'hbb2c34bf),
	.w4(32'hbb065625),
	.w5(32'h3b18f901),
	.w6(32'hbb87c28b),
	.w7(32'hbb917b6f),
	.w8(32'hbc3d299b),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5949e5),
	.w1(32'h3ad5e351),
	.w2(32'h3bb64ffe),
	.w3(32'h399e038a),
	.w4(32'h381c32aa),
	.w5(32'hbaa12e99),
	.w6(32'hbc1e9cdd),
	.w7(32'hbba4df1d),
	.w8(32'hbb0d26b5),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b49d659),
	.w1(32'hbad61eba),
	.w2(32'h3aa7d0fc),
	.w3(32'hbb083751),
	.w4(32'h3be5b555),
	.w5(32'h3a6ebaf9),
	.w6(32'hbb83887b),
	.w7(32'hba90ecf7),
	.w8(32'hbbee4756),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0de8da),
	.w1(32'hbb292156),
	.w2(32'h3aa7facb),
	.w3(32'hb986b3bc),
	.w4(32'h3b1c1523),
	.w5(32'hba4277ea),
	.w6(32'hbbe9eafb),
	.w7(32'hbb32ac74),
	.w8(32'h3b09e338),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3383dd),
	.w1(32'h3c808fa2),
	.w2(32'h3c38d1cd),
	.w3(32'hbb57bc64),
	.w4(32'h3afc5a23),
	.w5(32'h3b093f08),
	.w6(32'hba927092),
	.w7(32'hba9ac3d0),
	.w8(32'h3b4bd280),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b84dee9),
	.w1(32'h3b794d98),
	.w2(32'h39bbdb1b),
	.w3(32'h3b51c818),
	.w4(32'hba1c43b5),
	.w5(32'hba6e5c82),
	.w6(32'h3c1ef339),
	.w7(32'h3a9cd57c),
	.w8(32'hbb852e01),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb82b1da),
	.w1(32'hbaf71feb),
	.w2(32'hba9f8d7c),
	.w3(32'h3b2fac93),
	.w4(32'hbb2f203f),
	.w5(32'h3b598e67),
	.w6(32'h3b260819),
	.w7(32'h3a3ecd08),
	.w8(32'hbb8b4c44),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac7b5e4),
	.w1(32'hbbacfb62),
	.w2(32'hbb002c2f),
	.w3(32'hbbd7e97a),
	.w4(32'hbb2e5389),
	.w5(32'hbba177f2),
	.w6(32'hbbff1a43),
	.w7(32'hbbba3568),
	.w8(32'hbb4be891),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb32e184),
	.w1(32'hba3a5109),
	.w2(32'hba926fb9),
	.w3(32'hbae74022),
	.w4(32'hbbe56182),
	.w5(32'h3ba69fbc),
	.w6(32'h3aaae6c2),
	.w7(32'hbb8a00de),
	.w8(32'h3c3617d4),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2f2ce8),
	.w1(32'hbb0ae777),
	.w2(32'hbba3c055),
	.w3(32'h3c15a29d),
	.w4(32'hb8f17f94),
	.w5(32'h3b34f84f),
	.w6(32'h3b4c01ad),
	.w7(32'hbaf3b92a),
	.w8(32'h3ae0bf9c),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8410c8f),
	.w1(32'hba046a0e),
	.w2(32'h3a383605),
	.w3(32'h391b6768),
	.w4(32'h3a545f44),
	.w5(32'h3b4fee3a),
	.w6(32'h3a7c124b),
	.w7(32'hba0f38ac),
	.w8(32'hbbeb8402),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395776f4),
	.w1(32'hbb04b8e5),
	.w2(32'hbb8d7541),
	.w3(32'hba41ed9c),
	.w4(32'h3b265e8a),
	.w5(32'h3aa09a0d),
	.w6(32'hbc4bea5f),
	.w7(32'hbbe9d3a9),
	.w8(32'hb9c28f58),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b023cb0),
	.w1(32'h3b611ac3),
	.w2(32'h3b3f15b1),
	.w3(32'hb9abac5c),
	.w4(32'hba3a3cd4),
	.w5(32'hbab9fc38),
	.w6(32'h3b9fc097),
	.w7(32'h3ae866c8),
	.w8(32'hbb947662),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba830faf),
	.w1(32'h3a8e635b),
	.w2(32'h3b387dd0),
	.w3(32'hbafcb531),
	.w4(32'h3b0e60c0),
	.w5(32'hbb8929c8),
	.w6(32'h3ab68c5c),
	.w7(32'h3b3b6b79),
	.w8(32'hbae6b3dc),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9625bc),
	.w1(32'hbb3fe944),
	.w2(32'hbb7ae0c8),
	.w3(32'h3a6b5d73),
	.w4(32'hbb5cbc20),
	.w5(32'hbabc0fa1),
	.w6(32'h3a888726),
	.w7(32'hbab13b0c),
	.w8(32'hbb0da801),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a025e0d),
	.w1(32'h3b002b2e),
	.w2(32'h3b22f765),
	.w3(32'hbabd0ee5),
	.w4(32'h3a8810a3),
	.w5(32'h3b8e6f55),
	.w6(32'h3acf1532),
	.w7(32'h3b0f40bf),
	.w8(32'h3b496c75),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7c6fac),
	.w1(32'h3b428827),
	.w2(32'h3b35fe0c),
	.w3(32'h3ae1c7e4),
	.w4(32'hb9bfc60c),
	.w5(32'h3b1945dc),
	.w6(32'h3bc38374),
	.w7(32'h3adfca0a),
	.w8(32'hbb068469),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba926102),
	.w1(32'hb9278568),
	.w2(32'h3a607d5f),
	.w3(32'hba80bf02),
	.w4(32'h37a94c2b),
	.w5(32'h3c27e67b),
	.w6(32'h3abbcaea),
	.w7(32'h39d3c3c8),
	.w8(32'h3c57f5ec),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b62b3a7),
	.w1(32'h3be1005c),
	.w2(32'hb913db14),
	.w3(32'h3c5e3996),
	.w4(32'h3c181837),
	.w5(32'h3b90de6c),
	.w6(32'h3c8fc0bb),
	.w7(32'h3c129459),
	.w8(32'h39a8698d),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6ce1f72),
	.w1(32'h3a50fa09),
	.w2(32'h3bdfd3d1),
	.w3(32'h3a380437),
	.w4(32'h3c011ca6),
	.w5(32'h391f9b4d),
	.w6(32'hbbaacf32),
	.w7(32'h3abffbf1),
	.w8(32'hba6950b4),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a708393),
	.w1(32'hbac77121),
	.w2(32'hbb819bd3),
	.w3(32'hbb2645d1),
	.w4(32'h3a39acd1),
	.w5(32'hb88e57f8),
	.w6(32'hbc0b7da9),
	.w7(32'hbb3d2fe1),
	.w8(32'hba4959f2),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb542ab6),
	.w1(32'hbacab225),
	.w2(32'hbb000d25),
	.w3(32'h3aefe821),
	.w4(32'hba942648),
	.w5(32'h39c5ac25),
	.w6(32'h3b8674b1),
	.w7(32'hbac3c492),
	.w8(32'h3b112d6c),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8fb05d),
	.w1(32'h3a94316f),
	.w2(32'hbb8336d9),
	.w3(32'h3a40bc59),
	.w4(32'hbabf4349),
	.w5(32'h3b8e467c),
	.w6(32'h3b4ee345),
	.w7(32'hba83bc87),
	.w8(32'h3b894403),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2f4e4f),
	.w1(32'h3b1008b8),
	.w2(32'h3b66442f),
	.w3(32'h3c197098),
	.w4(32'h3bc9a041),
	.w5(32'hb96567b2),
	.w6(32'h3c77e99f),
	.w7(32'h3bfb7104),
	.w8(32'hbb351db9),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6caa35),
	.w1(32'hbbb18202),
	.w2(32'hbb90bc49),
	.w3(32'hbb96a903),
	.w4(32'hbb67ba29),
	.w5(32'h3b9ecf95),
	.w6(32'hbb2949da),
	.w7(32'hbbb0d0da),
	.w8(32'h3b639c63),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaef2947),
	.w1(32'hb9cc8aaf),
	.w2(32'h39ce06e8),
	.w3(32'h39ce0309),
	.w4(32'hbb980250),
	.w5(32'h3afb2be4),
	.w6(32'hbb004aa0),
	.w7(32'hbadfaa39),
	.w8(32'h3ba0baef),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2e7a9f),
	.w1(32'h3ba3ab94),
	.w2(32'h3934e0ed),
	.w3(32'hbb5411b2),
	.w4(32'h3a90e180),
	.w5(32'h39ec286f),
	.w6(32'hbc0ddd42),
	.w7(32'hba9c7fa0),
	.w8(32'h3aeb2747),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b978747),
	.w1(32'h3b00894c),
	.w2(32'h3a9858cc),
	.w3(32'hba8965ca),
	.w4(32'h3a53e14d),
	.w5(32'h3b697776),
	.w6(32'hbad08331),
	.w7(32'h3b0e8366),
	.w8(32'h3b8727dc),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbed1ae),
	.w1(32'h3b9143d7),
	.w2(32'h3bf48dfb),
	.w3(32'h399e93c6),
	.w4(32'h3b9b52a7),
	.w5(32'h39f9d2e0),
	.w6(32'h3b7149d7),
	.w7(32'h3bb7483c),
	.w8(32'hbc1b99d3),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adda3d2),
	.w1(32'hbb28c44a),
	.w2(32'h3ae869fe),
	.w3(32'hbc1c5aa1),
	.w4(32'hbbd5cbb7),
	.w5(32'hbb8021c5),
	.w6(32'hbc8b8d14),
	.w7(32'hbc1d4333),
	.w8(32'hbb80e90d),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaef2533),
	.w1(32'h3a15462f),
	.w2(32'h3b6a99d8),
	.w3(32'hbb8da156),
	.w4(32'h3b1d0de4),
	.w5(32'h3c06b5cf),
	.w6(32'hbbc079b0),
	.w7(32'h3ab1f100),
	.w8(32'h3c246344),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aef1ea6),
	.w1(32'h3b7c749e),
	.w2(32'h3b092cf8),
	.w3(32'h3c66cb7e),
	.w4(32'h3b03009d),
	.w5(32'h39ff7505),
	.w6(32'h3c2e19d8),
	.w7(32'h3af1fee8),
	.w8(32'h3b82b523),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad5c698),
	.w1(32'h3b9948d3),
	.w2(32'h3a043f02),
	.w3(32'h3bb11945),
	.w4(32'h3a5a6ff9),
	.w5(32'h3aefabd4),
	.w6(32'h3c9aa84f),
	.w7(32'h3bebaa05),
	.w8(32'h3b92b8c4),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5c0c42),
	.w1(32'hbb3da468),
	.w2(32'hbb2bf443),
	.w3(32'hba139e7a),
	.w4(32'h3b72b3b1),
	.w5(32'hbb869f60),
	.w6(32'h3bc01548),
	.w7(32'h3b646e77),
	.w8(32'hbbf96e9d),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5a836a),
	.w1(32'hbbab42c7),
	.w2(32'hbbea6294),
	.w3(32'hbbeda6dc),
	.w4(32'hbbc3a6d1),
	.w5(32'h3c11c427),
	.w6(32'hbbe10212),
	.w7(32'hbc09c6cb),
	.w8(32'h3c6461b9),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c710e79),
	.w1(32'h3c8af588),
	.w2(32'h3af04508),
	.w3(32'h3b1f2232),
	.w4(32'h3b94987f),
	.w5(32'h39d66a3b),
	.w6(32'h3b910746),
	.w7(32'hbb3ad9f2),
	.w8(32'h3b13a4c1),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b244350),
	.w1(32'hbaa34628),
	.w2(32'hba99f1a0),
	.w3(32'hbb80ac6c),
	.w4(32'h3ac79e65),
	.w5(32'hbbac9f8d),
	.w6(32'hbbbb571b),
	.w7(32'h3a7d03a1),
	.w8(32'h3aebfe89),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c48cd28),
	.w1(32'h3c850168),
	.w2(32'h3c297686),
	.w3(32'hbb8a587b),
	.w4(32'hba951662),
	.w5(32'h3c76761c),
	.w6(32'h394a6a76),
	.w7(32'h3a5431e6),
	.w8(32'h3c804fdc),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdcc2fb),
	.w1(32'hba0174c1),
	.w2(32'h3aff9c2f),
	.w3(32'h3cc3f33f),
	.w4(32'h3c7c9ba4),
	.w5(32'hb9f4169c),
	.w6(32'h3c8b0972),
	.w7(32'h3c22b7b4),
	.w8(32'hba2f7a14),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af5cb9a),
	.w1(32'h3c07ebc1),
	.w2(32'h3b875557),
	.w3(32'h3c17cd8e),
	.w4(32'h3b21c0ce),
	.w5(32'h3a148407),
	.w6(32'h3bba6625),
	.w7(32'h3bfbadb4),
	.w8(32'hbba16255),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb11fd3f),
	.w1(32'hbb5b4e18),
	.w2(32'hbacfd72b),
	.w3(32'hbb2c5824),
	.w4(32'hb91e125c),
	.w5(32'h3ca1dfa3),
	.w6(32'hbb4a8ca8),
	.w7(32'h38b77d61),
	.w8(32'h3b633d22),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b381c07),
	.w1(32'hbb5790f2),
	.w2(32'hba360bd9),
	.w3(32'h3c9a9777),
	.w4(32'h3c21ebe2),
	.w5(32'h3b224d53),
	.w6(32'h3b5fce59),
	.w7(32'h3c1ef0b3),
	.w8(32'h3a985537),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad0ab0f),
	.w1(32'h3b99f997),
	.w2(32'h3c3efd3d),
	.w3(32'h3b31bc34),
	.w4(32'h3bbfeaf7),
	.w5(32'hba37db76),
	.w6(32'h3b7785f9),
	.w7(32'h3c1223ab),
	.w8(32'h3b830fe3),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf48a38),
	.w1(32'h3c5c592b),
	.w2(32'h3bc61b32),
	.w3(32'hb8976009),
	.w4(32'h3af33fbd),
	.w5(32'h3ae0ec4d),
	.w6(32'h3bc6f402),
	.w7(32'hba9be2dd),
	.w8(32'h3b31b3cf),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b986626),
	.w1(32'h3b80c566),
	.w2(32'h3b904609),
	.w3(32'hbb441268),
	.w4(32'h3a81ca66),
	.w5(32'hbb09ddfc),
	.w6(32'h3a86e780),
	.w7(32'h3b3e40da),
	.w8(32'hbabc70bf),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb6cca4),
	.w1(32'hbab7714f),
	.w2(32'h3b0bdae8),
	.w3(32'hba477975),
	.w4(32'h3b237717),
	.w5(32'h3afd30aa),
	.w6(32'hbb2b350a),
	.w7(32'hbb0bf966),
	.w8(32'hba93ac4b),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2393ee),
	.w1(32'hbbc5fe65),
	.w2(32'hb9bc27af),
	.w3(32'hbb2c3f4b),
	.w4(32'hb90185c7),
	.w5(32'h3c1bd9ca),
	.w6(32'hbb88efec),
	.w7(32'hbb1984ad),
	.w8(32'h3bfeb32b),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bba3da5),
	.w1(32'h3bd9dc2b),
	.w2(32'h3ba31b48),
	.w3(32'h3ba9f9f3),
	.w4(32'hba02de74),
	.w5(32'h3b6812df),
	.w6(32'h3c00d60d),
	.w7(32'h3bb8e950),
	.w8(32'h3bee329e),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf28c20),
	.w1(32'h3b6f6c0c),
	.w2(32'hbabadfb8),
	.w3(32'h3bea3c49),
	.w4(32'hb9d4f238),
	.w5(32'h3b2c8886),
	.w6(32'h3ca00dca),
	.w7(32'h3bac72fd),
	.w8(32'hbb1191a1),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb19ec5e),
	.w1(32'hbb051272),
	.w2(32'hbb1969f9),
	.w3(32'h3b3cdd0b),
	.w4(32'h3b829cf9),
	.w5(32'hbb27c3b5),
	.w6(32'hbb95c345),
	.w7(32'hbb96b357),
	.w8(32'h3a9821e7),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb22a683),
	.w1(32'h3b2fb5ba),
	.w2(32'hbbabc608),
	.w3(32'h3b65ecf0),
	.w4(32'hbb4e7add),
	.w5(32'hbb456258),
	.w6(32'h3c5507a7),
	.w7(32'h3ae11c42),
	.w8(32'h3bff1ba4),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba74ee40),
	.w1(32'h3c1bf276),
	.w2(32'hba6dcc83),
	.w3(32'h3b8e830a),
	.w4(32'hbbdc3542),
	.w5(32'h3bfec9d5),
	.w6(32'h3cbae826),
	.w7(32'h3bd76265),
	.w8(32'h3c2010b6),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c10ffd9),
	.w1(32'h3c10b2a2),
	.w2(32'h3bac07e0),
	.w3(32'h3bf57451),
	.w4(32'h3b84f4e4),
	.w5(32'h3ba2aad8),
	.w6(32'h3c89c725),
	.w7(32'h3c21b3c3),
	.w8(32'h3c442efa),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b66104d),
	.w1(32'h3b846feb),
	.w2(32'hbaaf3917),
	.w3(32'h3af617dc),
	.w4(32'hbb1f8c40),
	.w5(32'h3b821d00),
	.w6(32'h3c57e725),
	.w7(32'h3bb339fc),
	.w8(32'h3ac67993),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba9e47a),
	.w1(32'h3b8acff7),
	.w2(32'h3bd917c6),
	.w3(32'h3b41e73f),
	.w4(32'h3b953e27),
	.w5(32'hbae1f488),
	.w6(32'h3a4ed2cc),
	.w7(32'h3b1b6eb5),
	.w8(32'hbba4eea4),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb982e7ba),
	.w1(32'hbb109aa4),
	.w2(32'h3470e726),
	.w3(32'hbbb2d83a),
	.w4(32'hbb38e899),
	.w5(32'h3b5e1467),
	.w6(32'hbc00477a),
	.w7(32'hbbd738b8),
	.w8(32'h3b12a3a0),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38085497),
	.w1(32'hbb43b08a),
	.w2(32'h3a708da2),
	.w3(32'hbab50b31),
	.w4(32'h3ae01592),
	.w5(32'hbc8a3c4a),
	.w6(32'hb9ab7ce3),
	.w7(32'h3ac37d5f),
	.w8(32'hbc17167b),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3dc2a2),
	.w1(32'hba8b9338),
	.w2(32'hbb4f89e5),
	.w3(32'hbb8294ff),
	.w4(32'hbbaddcea),
	.w5(32'hbbb752cf),
	.w6(32'hbb97b7ec),
	.w7(32'hbb10479f),
	.w8(32'hbb1d5bbc),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2f0e3c),
	.w1(32'hba65f0a1),
	.w2(32'hbb93d606),
	.w3(32'hbc121411),
	.w4(32'hbbef4fcb),
	.w5(32'h3bdd4415),
	.w6(32'hbbcecab3),
	.w7(32'hbbaf03f4),
	.w8(32'h3c504bbd),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb285090),
	.w1(32'h3b910e6d),
	.w2(32'h3a8c8056),
	.w3(32'h3c904f47),
	.w4(32'h39738e2a),
	.w5(32'h3b7476be),
	.w6(32'h3ca628f0),
	.w7(32'h3b3251d1),
	.w8(32'h3b0d8d65),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6fbddf),
	.w1(32'h3c0067c7),
	.w2(32'h3b2d8646),
	.w3(32'h3b034a56),
	.w4(32'h3b48989d),
	.w5(32'h3bb5546a),
	.w6(32'h3c208a35),
	.w7(32'hb9d312f3),
	.w8(32'h3bcdf9c1),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b806590),
	.w1(32'h3b8de378),
	.w2(32'hb9c6b4fc),
	.w3(32'h3c248661),
	.w4(32'h3c29208f),
	.w5(32'h3a207f32),
	.w6(32'h3ba5926c),
	.w7(32'h3c4ccdf9),
	.w8(32'h3a8c4038),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb88dedf),
	.w1(32'hbba80db6),
	.w2(32'hbb33fe1d),
	.w3(32'h37e9d8aa),
	.w4(32'h3a5f20aa),
	.w5(32'h3c3e241f),
	.w6(32'h3b9a0a38),
	.w7(32'h3baa17b6),
	.w8(32'h3c29f482),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c165bc7),
	.w1(32'h3c0ed53a),
	.w2(32'h3c32c173),
	.w3(32'h3c089391),
	.w4(32'h3c17d812),
	.w5(32'h3c0c1398),
	.w6(32'h3c7628df),
	.w7(32'h3c921768),
	.w8(32'h3c5ef6ff),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bff6c0c),
	.w1(32'h3b95b52d),
	.w2(32'hbb39f9fa),
	.w3(32'h3ab9ecc5),
	.w4(32'hbb3c9357),
	.w5(32'hba62863f),
	.w6(32'hbb543214),
	.w7(32'hbba9f00d),
	.w8(32'hbb24e1f6),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb70890d),
	.w1(32'hbb98fccb),
	.w2(32'hba4e33ed),
	.w3(32'hbb99cb7e),
	.w4(32'h3a06186b),
	.w5(32'h3b0e24ab),
	.w6(32'hbac0d2da),
	.w7(32'h3a293fcc),
	.w8(32'h3c05332b),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbfc072),
	.w1(32'h3c4581cc),
	.w2(32'h3c0149f4),
	.w3(32'h3b2752c2),
	.w4(32'h3a99d6df),
	.w5(32'hba23c339),
	.w6(32'h3c19a0b3),
	.w7(32'h3c2d4dcc),
	.w8(32'h390e5452),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba2c7de),
	.w1(32'hbae9c517),
	.w2(32'hbb45fa65),
	.w3(32'h389edd0e),
	.w4(32'h3ab72c8e),
	.w5(32'h3b83a289),
	.w6(32'hba9c4eea),
	.w7(32'hbb1ebb1b),
	.w8(32'h3b82d129),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9b0287),
	.w1(32'h3b9001a4),
	.w2(32'hba4d6988),
	.w3(32'h3bde8b3a),
	.w4(32'h3aa819b1),
	.w5(32'h3b20ff84),
	.w6(32'h3c5503a7),
	.w7(32'h3b297fde),
	.w8(32'h3c02627b),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a29a5bf),
	.w1(32'hbb08787b),
	.w2(32'hbbd2f0c8),
	.w3(32'h3b816d83),
	.w4(32'hbbab5324),
	.w5(32'hbb408c37),
	.w6(32'h3be9c5b1),
	.w7(32'h3b9b5e7a),
	.w8(32'hbbc616d1),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d4877),
	.w1(32'hbba0c74a),
	.w2(32'hbb94f25b),
	.w3(32'hbba14e0e),
	.w4(32'hbbc99f08),
	.w5(32'h3b9ce6d5),
	.w6(32'hbb9cfbca),
	.w7(32'hbabbdbeb),
	.w8(32'h3b08b9eb),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4da928),
	.w1(32'hb9bb60f7),
	.w2(32'h3b173cad),
	.w3(32'h3bbdd824),
	.w4(32'h3c101cf6),
	.w5(32'h3c16e368),
	.w6(32'h3ab7ceb0),
	.w7(32'h3ca3d326),
	.w8(32'h3c0bf019),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b19da5d),
	.w1(32'h3bdcfb54),
	.w2(32'h39909149),
	.w3(32'h3c824748),
	.w4(32'h3b8158db),
	.w5(32'h3bd62a14),
	.w6(32'h3c5e8ff5),
	.w7(32'h3bdcb86a),
	.w8(32'h3be0033f),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8d807e),
	.w1(32'hbb5b79f2),
	.w2(32'hbbc8140d),
	.w3(32'h3bc23a1b),
	.w4(32'hb84c3a1e),
	.w5(32'hbc52c156),
	.w6(32'h3b4fb028),
	.w7(32'hbb1c6d27),
	.w8(32'hbbd4190b),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf26b7e),
	.w1(32'h381fc0c3),
	.w2(32'h3b1f8745),
	.w3(32'hbb923fb5),
	.w4(32'hb9f6a4f9),
	.w5(32'hba20165a),
	.w6(32'h3bb548db),
	.w7(32'h3b963d6c),
	.w8(32'hbb364bd6),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae3d5e6),
	.w1(32'h38e61ad5),
	.w2(32'h3b419a88),
	.w3(32'h3bc19fd2),
	.w4(32'h3c19ae83),
	.w5(32'hba23ba38),
	.w6(32'h3a23a017),
	.w7(32'h3cb2c3b0),
	.w8(32'hbbe75d27),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9e4930),
	.w1(32'hbbe0f741),
	.w2(32'h3b0e215d),
	.w3(32'hbb8cd627),
	.w4(32'h3996e025),
	.w5(32'h3b1cbf5a),
	.w6(32'hbb4682a7),
	.w7(32'hba815573),
	.w8(32'hb81692c8),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a929022),
	.w1(32'h3b75943e),
	.w2(32'h3af65550),
	.w3(32'h3b57ce5b),
	.w4(32'h3ba47b9d),
	.w5(32'h3b89d341),
	.w6(32'h3b1f7798),
	.w7(32'h3931500c),
	.w8(32'hba556ff5),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa08f7d),
	.w1(32'hbb350bf7),
	.w2(32'hbba4e217),
	.w3(32'h3b8e8778),
	.w4(32'hb7984980),
	.w5(32'h3b382435),
	.w6(32'h3a7b10b5),
	.w7(32'h3a66afe6),
	.w8(32'hbbb59f50),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390be694),
	.w1(32'hbb248fdf),
	.w2(32'h37853d57),
	.w3(32'h3b069982),
	.w4(32'h3b1fc8fc),
	.w5(32'hbb1c7470),
	.w6(32'hbbc167ab),
	.w7(32'hbb1ed7d7),
	.w8(32'hbb49d053),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2675fa),
	.w1(32'hbb2f4d2b),
	.w2(32'hbb60384f),
	.w3(32'hbbf487d3),
	.w4(32'hbba45e91),
	.w5(32'h3c3fb193),
	.w6(32'hbbf8c643),
	.w7(32'hbb9d9897),
	.w8(32'h3c292ea6),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bde0dd1),
	.w1(32'h39ef2bdf),
	.w2(32'h3a6b24c4),
	.w3(32'h3bb202ed),
	.w4(32'h3b493f48),
	.w5(32'h3ba493b5),
	.w6(32'h3b9d870f),
	.w7(32'h3a285d9a),
	.w8(32'hbb228ee1),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af62f2e),
	.w1(32'h3b1e9616),
	.w2(32'h3b602c36),
	.w3(32'h3a185593),
	.w4(32'h3b693272),
	.w5(32'h3b98e360),
	.w6(32'hbbcd6dc3),
	.w7(32'hbb31a5e4),
	.w8(32'hba88edf4),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0cbee6),
	.w1(32'h3c322752),
	.w2(32'h3c0fb5d2),
	.w3(32'hbad8faf3),
	.w4(32'hbae7e8fd),
	.w5(32'hbc0846c9),
	.w6(32'hbbac38ab),
	.w7(32'hba82aa82),
	.w8(32'hbbcace56),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfa3f0a),
	.w1(32'hbbd294dc),
	.w2(32'hbc05bb53),
	.w3(32'hbbb2cd4e),
	.w4(32'hbb80650a),
	.w5(32'h3ba26ed6),
	.w6(32'hbadcef0d),
	.w7(32'hbad039d4),
	.w8(32'h3a895536),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afc1328),
	.w1(32'hba3d0b3e),
	.w2(32'h3ae09616),
	.w3(32'h38b751e2),
	.w4(32'hba8a04bd),
	.w5(32'h3bbaa864),
	.w6(32'hbaff9f70),
	.w7(32'hb9392840),
	.w8(32'h3b667258),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf15b03),
	.w1(32'h3c04efc2),
	.w2(32'h3be77da5),
	.w3(32'h3be34b1d),
	.w4(32'h3b87faa3),
	.w5(32'h3b2e380c),
	.w6(32'h3c249820),
	.w7(32'h3b7e8549),
	.w8(32'hbaa7080a),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b15feac),
	.w1(32'h3b0a0b22),
	.w2(32'h3ba8e12d),
	.w3(32'h3b3b6cf7),
	.w4(32'h3bb21d91),
	.w5(32'h3b14a10a),
	.w6(32'hbc03ef7d),
	.w7(32'h3aa34e23),
	.w8(32'hbb81955a),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2f1ddb),
	.w1(32'hbb3c236b),
	.w2(32'h3b354d6e),
	.w3(32'h3a07551f),
	.w4(32'h3a773715),
	.w5(32'h3bf6799e),
	.w6(32'hbb9df0cc),
	.w7(32'hbb60fd2b),
	.w8(32'hbb9f09b3),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd1c496),
	.w1(32'h3c060438),
	.w2(32'h3c6c2238),
	.w3(32'hbb4bc624),
	.w4(32'h3b77a14a),
	.w5(32'hbb26f79a),
	.w6(32'hbc05df13),
	.w7(32'h3c070c85),
	.w8(32'hba7c1ff3),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb78a4fa),
	.w1(32'h3a94b719),
	.w2(32'hba7e67dc),
	.w3(32'h3b20a03a),
	.w4(32'hbaaa26ae),
	.w5(32'h3bc05697),
	.w6(32'h3babc6de),
	.w7(32'h3af3e7a8),
	.w8(32'hbb82458e),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0f1d1a),
	.w1(32'h3b30746c),
	.w2(32'h3be9cd51),
	.w3(32'hbb43724b),
	.w4(32'hb9d7b019),
	.w5(32'h3bf0eb4d),
	.w6(32'hbc0a21e5),
	.w7(32'hbb8677e0),
	.w8(32'h3ae15cbd),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcd953b),
	.w1(32'h3bc66e2d),
	.w2(32'h3b6456cb),
	.w3(32'h3ba37d87),
	.w4(32'h3b3db308),
	.w5(32'h3b229cac),
	.w6(32'h3b7ac500),
	.w7(32'h3b17ef35),
	.w8(32'h3c0569c0),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a10fa51),
	.w1(32'h3b709a0e),
	.w2(32'hbb85d267),
	.w3(32'h3bbdeebb),
	.w4(32'h3b17f397),
	.w5(32'hbbeb807d),
	.w6(32'h3c61d351),
	.w7(32'h3b38a36b),
	.w8(32'h3b6a4d65),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4ec354),
	.w1(32'h3c2d0b44),
	.w2(32'h3b92ef57),
	.w3(32'hbc2bb794),
	.w4(32'hbc0208bf),
	.w5(32'h3b6ec2ab),
	.w6(32'hbb214b90),
	.w7(32'hbb995a8e),
	.w8(32'h3b2f7ff9),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8df119),
	.w1(32'h3b47e9f1),
	.w2(32'h399e9aa3),
	.w3(32'h3b8d2639),
	.w4(32'h3a54a4be),
	.w5(32'h3b34901e),
	.w6(32'h3c22016e),
	.w7(32'h3aa79f23),
	.w8(32'hba90c586),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7f6884),
	.w1(32'hbb5f15c4),
	.w2(32'h380248a8),
	.w3(32'hbb5e8168),
	.w4(32'hb8de0e49),
	.w5(32'hbb87018b),
	.w6(32'hbbebb028),
	.w7(32'hbace997d),
	.w8(32'hbba8f9fd),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3713dc58),
	.w1(32'h3a8f702d),
	.w2(32'h3ace56f5),
	.w3(32'hbaac480f),
	.w4(32'h3b0e4a34),
	.w5(32'h3bac3617),
	.w6(32'hbb843a03),
	.w7(32'hbb29ab84),
	.w8(32'h3bf4dfbd),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc6da5f),
	.w1(32'h3a81452d),
	.w2(32'hba376599),
	.w3(32'h3a7f9602),
	.w4(32'h3a4bbeb3),
	.w5(32'h3a88fa8a),
	.w6(32'hbb6299e5),
	.w7(32'h3ab3042d),
	.w8(32'h3ab2a456),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbde552d),
	.w1(32'hbb3cb3f6),
	.w2(32'hbb9755e4),
	.w3(32'h3bb94cde),
	.w4(32'h3b6c7266),
	.w5(32'h3c1744df),
	.w6(32'h3c4c0744),
	.w7(32'h3bce37b5),
	.w8(32'h3c53900b),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acb6a0b),
	.w1(32'h3ab1a606),
	.w2(32'hbc25f676),
	.w3(32'h3c47764b),
	.w4(32'hbb051cde),
	.w5(32'h3b8b86d5),
	.w6(32'h3c16583e),
	.w7(32'hbb333c10),
	.w8(32'h3ba8dcf3),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbc880c),
	.w1(32'h3b3c8d98),
	.w2(32'h3abdf313),
	.w3(32'h3b8fb559),
	.w4(32'h3b32897f),
	.w5(32'h3b2b8014),
	.w6(32'h3b4fee33),
	.w7(32'h3b4c116f),
	.w8(32'h3be91ba8),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf6441d),
	.w1(32'hbb57b35e),
	.w2(32'h3b0495c5),
	.w3(32'h3b8b96ec),
	.w4(32'h3bc20b05),
	.w5(32'h3b4ba8a4),
	.w6(32'h3b93fed2),
	.w7(32'h3b7e0387),
	.w8(32'h3ab0c26e),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1d279c),
	.w1(32'h3ae612f3),
	.w2(32'h3b0ebd57),
	.w3(32'hbad7c19f),
	.w4(32'hbac40a83),
	.w5(32'hbbdabde2),
	.w6(32'hbb06db5a),
	.w7(32'h38296b2a),
	.w8(32'hbbbaf71f),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9e0748),
	.w1(32'h3c3e27a5),
	.w2(32'h3b978b3a),
	.w3(32'h3ad5f258),
	.w4(32'hbb4317ac),
	.w5(32'h3ad30e9e),
	.w6(32'h38e94e74),
	.w7(32'h3bdbd20d),
	.w8(32'h3b902709),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b812fbe),
	.w1(32'hbb9183d5),
	.w2(32'hbb49a414),
	.w3(32'hbb955305),
	.w4(32'hbb4fd8fe),
	.w5(32'h3b3376f3),
	.w6(32'hba9c217b),
	.w7(32'hbb092f29),
	.w8(32'h3b8495f7),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7d2bfb),
	.w1(32'h3b44eba8),
	.w2(32'hb9981b92),
	.w3(32'h3b2e4ec2),
	.w4(32'hbbaf6ebe),
	.w5(32'hbc2f4078),
	.w6(32'h3c05bbec),
	.w7(32'h3b35b858),
	.w8(32'hbb87068a),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd93809),
	.w1(32'hbb85042a),
	.w2(32'hbc18354e),
	.w3(32'hbc038e41),
	.w4(32'hbc1e0234),
	.w5(32'h3ac1ca3e),
	.w6(32'h3bca4432),
	.w7(32'hbb563b57),
	.w8(32'hbb6f245d),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0347c9),
	.w1(32'h3beab201),
	.w2(32'h3bb62acb),
	.w3(32'hbb9b8770),
	.w4(32'hbbc5721a),
	.w5(32'h3b8fbb54),
	.w6(32'hbbeb2190),
	.w7(32'hbb26b16c),
	.w8(32'h3b8b00fe),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4315ca),
	.w1(32'hbb9ccbf6),
	.w2(32'h3af2834f),
	.w3(32'hbadf8155),
	.w4(32'h3ab26ff4),
	.w5(32'hbca4c394),
	.w6(32'hbbc81afa),
	.w7(32'h3b1ca5f7),
	.w8(32'hbc543a3c),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc918384),
	.w1(32'hbc45fde4),
	.w2(32'hbc8961f0),
	.w3(32'hbc4bcc37),
	.w4(32'hbcb7c420),
	.w5(32'hbb94fc31),
	.w6(32'hbb762a88),
	.w7(32'hbc62d9dd),
	.w8(32'h3ba2cbfc),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b7351),
	.w1(32'hbb8f6461),
	.w2(32'hbb2617dd),
	.w3(32'hbc5d48a1),
	.w4(32'hbc416e83),
	.w5(32'hbbb7fde2),
	.w6(32'hb99f6533),
	.w7(32'hbc0ec988),
	.w8(32'hbb34fb1a),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb34cd4a),
	.w1(32'hbb5734dd),
	.w2(32'hbb37a607),
	.w3(32'hbad2f980),
	.w4(32'h3a3b1cc4),
	.w5(32'hb9bd913f),
	.w6(32'hba9cfe1c),
	.w7(32'h3a701495),
	.w8(32'h3c064c00),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af33ce8),
	.w1(32'hbac8abf5),
	.w2(32'hbc28bd65),
	.w3(32'hbb382d7e),
	.w4(32'hbb89e104),
	.w5(32'h39499c44),
	.w6(32'h3bbd363c),
	.w7(32'hbb68c8ae),
	.w8(32'hbb4c7329),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae2bc38),
	.w1(32'hbb4a5d14),
	.w2(32'h3b02b66d),
	.w3(32'hbb48e83f),
	.w4(32'hbaab64c5),
	.w5(32'h3c5472bd),
	.w6(32'hbc27cc2e),
	.w7(32'h39807375),
	.w8(32'h3c78407e),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c830d15),
	.w1(32'h3c1a1401),
	.w2(32'hbbdcfd16),
	.w3(32'h3c237e17),
	.w4(32'hbb9f5c65),
	.w5(32'h3c01189e),
	.w6(32'h3c550658),
	.w7(32'hbba7119d),
	.w8(32'hbc00ce0b),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0f3b9e),
	.w1(32'hbcafcfcf),
	.w2(32'h3a8ef339),
	.w3(32'hbc70f420),
	.w4(32'h3ba94088),
	.w5(32'hbb15dc82),
	.w6(32'hbd2625dc),
	.w7(32'hbc7726ac),
	.w8(32'hbbba01a1),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8e4a8c),
	.w1(32'hbc2e5ae7),
	.w2(32'hbc060020),
	.w3(32'hbc1436b5),
	.w4(32'hbbb2bce7),
	.w5(32'h3bca9397),
	.w6(32'hbc8cee1e),
	.w7(32'hbc2e5a5c),
	.w8(32'h3a34d640),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8cfa54),
	.w1(32'hbaf70147),
	.w2(32'h3aff5edb),
	.w3(32'h3b2319f7),
	.w4(32'hbb5725a5),
	.w5(32'h3ca57c5f),
	.w6(32'h39abcf5f),
	.w7(32'hb87b4c85),
	.w8(32'h3c2105bd),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c890bc4),
	.w1(32'h3b8d7db4),
	.w2(32'h3c9e1633),
	.w3(32'h3bae7521),
	.w4(32'h3ce7b5c4),
	.w5(32'h3b1ba810),
	.w6(32'hbc78a2d0),
	.w7(32'h3c6b02f3),
	.w8(32'h3b90880e),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a7b18f),
	.w1(32'hbb4a332f),
	.w2(32'h3b369b9a),
	.w3(32'hba3b0a41),
	.w4(32'h396d1c95),
	.w5(32'hbb955607),
	.w6(32'hba089420),
	.w7(32'hba56ffbf),
	.w8(32'hbbb6fca9),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5d2b52),
	.w1(32'hbb558e38),
	.w2(32'hbbe3d9c7),
	.w3(32'h3a8fbd34),
	.w4(32'hbc5d0ba3),
	.w5(32'h3b4b67bf),
	.w6(32'h38142936),
	.w7(32'h3adbdb85),
	.w8(32'hb9b09b16),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5c7cf7),
	.w1(32'hba6a62e8),
	.w2(32'h3b9a4177),
	.w3(32'hbaf974c4),
	.w4(32'hbb0e83ac),
	.w5(32'h3c43a0c4),
	.w6(32'hbb3c3151),
	.w7(32'hba9d5eb2),
	.w8(32'h3c1376c8),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6879c3),
	.w1(32'hba6271f1),
	.w2(32'h3a4694ec),
	.w3(32'h3c14760f),
	.w4(32'h3bf5a7e1),
	.w5(32'hbbfcf0ae),
	.w6(32'h3c050b91),
	.w7(32'h3acd5e1b),
	.w8(32'h3b5972d9),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb88f92a),
	.w1(32'h3ba61f11),
	.w2(32'hbb9aaed4),
	.w3(32'hbbbd3fce),
	.w4(32'hbb70910c),
	.w5(32'hbc4c7851),
	.w6(32'h3a7aaa9d),
	.w7(32'hbbe0211c),
	.w8(32'hbbe01df6),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc47a089),
	.w1(32'hbc894ffd),
	.w2(32'hbc50330e),
	.w3(32'hbc469007),
	.w4(32'hbc06af2e),
	.w5(32'h3bc98747),
	.w6(32'hbc2627a4),
	.w7(32'hbbd3256a),
	.w8(32'h3cc83afd),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb6d240),
	.w1(32'h3cdcaa69),
	.w2(32'h3b10884f),
	.w3(32'h3c865ab6),
	.w4(32'hb9afeffa),
	.w5(32'h3bda64f8),
	.w6(32'h3d2c79c3),
	.w7(32'h3c49cec0),
	.w8(32'h3aaa39ee),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96c03a6),
	.w1(32'hbb2b01bd),
	.w2(32'hbbd2e549),
	.w3(32'h3bb07a49),
	.w4(32'hbc0f2929),
	.w5(32'hbb03c44c),
	.w6(32'h392ad16b),
	.w7(32'hbc169c5f),
	.w8(32'hb9c2e3d6),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb3a346),
	.w1(32'h3b800f08),
	.w2(32'h3b9af809),
	.w3(32'h3afb9173),
	.w4(32'h37dd7900),
	.w5(32'hbae17f54),
	.w6(32'h3b6ed54c),
	.w7(32'h3b12652f),
	.w8(32'hbbfd308c),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393f4f0b),
	.w1(32'h3b41dafd),
	.w2(32'h37e83b5e),
	.w3(32'h3b9dfc64),
	.w4(32'h3bfd434f),
	.w5(32'h3b4d9cfc),
	.w6(32'hbc91ab71),
	.w7(32'hbb8e9c16),
	.w8(32'h39deb0a8),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b849e9a),
	.w1(32'hbadda0fa),
	.w2(32'h3b5e73a6),
	.w3(32'hba4e997c),
	.w4(32'h3b0678a6),
	.w5(32'hb9c5e57b),
	.w6(32'hbc7d7e36),
	.w7(32'h3b037a00),
	.w8(32'hbbfeff86),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb11b503),
	.w1(32'hbba9149d),
	.w2(32'hba21a6a5),
	.w3(32'h3a4dd022),
	.w4(32'h3bfe82ce),
	.w5(32'h3aa3437f),
	.w6(32'hbcaf5732),
	.w7(32'hbad6466d),
	.w8(32'hbb1f0299),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a811c54),
	.w1(32'hba0e5cc1),
	.w2(32'h3ba1f732),
	.w3(32'h3b2e79d0),
	.w4(32'h3ab4fa3a),
	.w5(32'h3acba476),
	.w6(32'hbbfe6d4e),
	.w7(32'h3a6682fb),
	.w8(32'hbb4ae7dd),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc0d046),
	.w1(32'hbb8ab218),
	.w2(32'h3a218ea6),
	.w3(32'hbb108d54),
	.w4(32'h3b7b8c16),
	.w5(32'hbb53c698),
	.w6(32'hbc8f35d6),
	.w7(32'hbb96192f),
	.w8(32'hbc07961e),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd14cd0),
	.w1(32'hbb6b3d2d),
	.w2(32'hbb552933),
	.w3(32'hb91753c5),
	.w4(32'hbb9cc347),
	.w5(32'h3ccbedd3),
	.w6(32'h3af392c4),
	.w7(32'h3a97f4b6),
	.w8(32'h3c4687fa),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule