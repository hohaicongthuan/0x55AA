module layer_10_featuremap_153(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38736b4c),
	.w1(32'h381925d4),
	.w2(32'hb75b364e),
	.w3(32'h3869d77b),
	.w4(32'h37566173),
	.w5(32'hb741fd24),
	.w6(32'h382bc645),
	.w7(32'hb758aee6),
	.w8(32'h3626f89e),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9de125),
	.w1(32'hbbf920bb),
	.w2(32'hbb59c45f),
	.w3(32'hbae4c93a),
	.w4(32'hbc07ffb1),
	.w5(32'hbbc5c8a4),
	.w6(32'h3a4e1fbc),
	.w7(32'hbbdb5456),
	.w8(32'hbba6f77d),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3725063d),
	.w1(32'h37502542),
	.w2(32'h372cbbcc),
	.w3(32'h3682fb16),
	.w4(32'h37094ce4),
	.w5(32'h36823083),
	.w6(32'hb6881f7e),
	.w7(32'hb6ac981c),
	.w8(32'hb6a37c04),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a759ea4),
	.w1(32'h3b451da9),
	.w2(32'h3b4bad3e),
	.w3(32'h3a2a52cb),
	.w4(32'h3ac99167),
	.w5(32'h3b1ab8f9),
	.w6(32'h3a0f3a8e),
	.w7(32'h3a505c93),
	.w8(32'h39f67c9e),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a6d9f1),
	.w1(32'h396d7f1b),
	.w2(32'h39eff1a8),
	.w3(32'hb75b0318),
	.w4(32'h38b449d1),
	.w5(32'h399534a4),
	.w6(32'hb86209ed),
	.w7(32'hb7adfef0),
	.w8(32'h38dfa3cd),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3787776b),
	.w1(32'hb836b214),
	.w2(32'hb8443348),
	.w3(32'h38a25f7b),
	.w4(32'h37445f47),
	.w5(32'h364c83ff),
	.w6(32'h39040164),
	.w7(32'h38a4f2b5),
	.w8(32'h37846424),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8a39eb),
	.w1(32'h3c88a9e1),
	.w2(32'hbbd31d26),
	.w3(32'h3bbcd758),
	.w4(32'h3c0449f9),
	.w5(32'hbc02450c),
	.w6(32'h3bf07d1d),
	.w7(32'h3ba569ae),
	.w8(32'hbc64686d),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6acbc6),
	.w1(32'hbb4c5ff2),
	.w2(32'hbc42289b),
	.w3(32'hbbddfe5a),
	.w4(32'hbc6d2fc3),
	.w5(32'hbc3382b5),
	.w6(32'hbca55765),
	.w7(32'hbc40c639),
	.w8(32'hbcb307ce),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a295a4f),
	.w1(32'h396c29f3),
	.w2(32'h397029bf),
	.w3(32'h3a80057c),
	.w4(32'h39b2e738),
	.w5(32'h39acd2ba),
	.w6(32'h3a918ab0),
	.w7(32'h3a305714),
	.w8(32'h385bf5e3),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1923b7),
	.w1(32'h3bfdaa9b),
	.w2(32'hbc2b258e),
	.w3(32'hb8619c22),
	.w4(32'h3bb75f1c),
	.w5(32'hbbf085f4),
	.w6(32'h3a90b950),
	.w7(32'h3b5b53b7),
	.w8(32'hbbfc68a4),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e9daee),
	.w1(32'h39f143f4),
	.w2(32'h39b92583),
	.w3(32'h39ddd10f),
	.w4(32'h3a17fd46),
	.w5(32'h39a913b6),
	.w6(32'h39dd4df4),
	.w7(32'h3a318702),
	.w8(32'h397562a7),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c19c87c),
	.w1(32'h3cd9a42d),
	.w2(32'hbb7f232c),
	.w3(32'h3b7a2e86),
	.w4(32'h3c8fd2f5),
	.w5(32'hbbe5de97),
	.w6(32'h3b4b20cf),
	.w7(32'h3c577594),
	.w8(32'hbc7885a2),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b93be44),
	.w1(32'h3c22d0ce),
	.w2(32'hbbcaeb99),
	.w3(32'hba954fa9),
	.w4(32'h3bcedc2e),
	.w5(32'hbbe10dae),
	.w6(32'hbbbad7cc),
	.w7(32'h39d7393c),
	.w8(32'hbc0e0170),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be708c0),
	.w1(32'hb85d9ceb),
	.w2(32'hbb82ccec),
	.w3(32'h3ba37046),
	.w4(32'hbb007ba9),
	.w5(32'hbb905e9a),
	.w6(32'hb8b7bf7b),
	.w7(32'hbb504a56),
	.w8(32'hbb8c8bbb),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba5c1b8),
	.w1(32'hbb6c190f),
	.w2(32'hbb043516),
	.w3(32'hb8bb7bce),
	.w4(32'hbb237d7b),
	.w5(32'hbb1be89c),
	.w6(32'h3b607902),
	.w7(32'h38bb6ff4),
	.w8(32'hbb082c31),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac70d6e),
	.w1(32'hbb9b3adc),
	.w2(32'hbc45d6d8),
	.w3(32'hba60f86e),
	.w4(32'hbba3b538),
	.w5(32'hbc3beec6),
	.w6(32'hbb666bab),
	.w7(32'hbc562a05),
	.w8(32'hbc573917),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38748947),
	.w1(32'h38df7ebf),
	.w2(32'h3884429d),
	.w3(32'h39763e30),
	.w4(32'h38ea0d4c),
	.w5(32'hb8b49c5c),
	.w6(32'h39dd77a5),
	.w7(32'h395bffa0),
	.w8(32'h39294135),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7d6307),
	.w1(32'h3c342d98),
	.w2(32'hbc6ecb0f),
	.w3(32'h3a8fd64a),
	.w4(32'h3b192bf9),
	.w5(32'hbc8ef222),
	.w6(32'hbc3bbedb),
	.w7(32'hbc11fd76),
	.w8(32'hbc8bb596),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b910d58),
	.w1(32'h3be3de78),
	.w2(32'hbbc3be27),
	.w3(32'hbac87dce),
	.w4(32'h3b0500b0),
	.w5(32'hbbdc9a2f),
	.w6(32'hbb9ef314),
	.w7(32'hbb0eae8b),
	.w8(32'hbbfd21aa),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9561b1e),
	.w1(32'h37793b31),
	.w2(32'h39c15402),
	.w3(32'hb99aba20),
	.w4(32'h389d2115),
	.w5(32'h39b72a01),
	.w6(32'hb9783d49),
	.w7(32'hb966ab9a),
	.w8(32'hb638284f),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399241a1),
	.w1(32'h3a08562d),
	.w2(32'h398a65a3),
	.w3(32'h39209313),
	.w4(32'hb8982cce),
	.w5(32'h3777e576),
	.w6(32'h392b7217),
	.w7(32'hb8c57180),
	.w8(32'hb87d7bc0),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba586555),
	.w1(32'hba3b45a6),
	.w2(32'h3b167aa8),
	.w3(32'h3932e902),
	.w4(32'hba0da1ff),
	.w5(32'h3af07c5b),
	.w6(32'h3b469c04),
	.w7(32'h3ac22eb7),
	.w8(32'h3b031593),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a270ece),
	.w1(32'h3bf37578),
	.w2(32'hbc7e5d33),
	.w3(32'hbc2f0fee),
	.w4(32'h3c253872),
	.w5(32'hbc809071),
	.w6(32'hbc4e396a),
	.w7(32'h3a05e051),
	.w8(32'hbc4081f2),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9dfec6),
	.w1(32'hb8938e5b),
	.w2(32'hbb82a825),
	.w3(32'hbaef1f38),
	.w4(32'h3af9f1b6),
	.w5(32'hb9abaf80),
	.w6(32'h3a0c1548),
	.w7(32'h3b2aab85),
	.w8(32'h38e10a5c),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc32f4f5),
	.w1(32'hbbdb1543),
	.w2(32'h3ba2731c),
	.w3(32'hbbc7b8b5),
	.w4(32'hbc0fb210),
	.w5(32'hb897defd),
	.w6(32'h3c06af9b),
	.w7(32'hbb7211f1),
	.w8(32'h3a37fce1),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8147a90),
	.w1(32'h39b4d08f),
	.w2(32'hb89ee402),
	.w3(32'hb8d9616f),
	.w4(32'hb8087eb8),
	.w5(32'hba0afbe9),
	.w6(32'hb933ef5a),
	.w7(32'hb9aeede9),
	.w8(32'hba198f33),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6c3eaea),
	.w1(32'h3809daa8),
	.w2(32'h3967a246),
	.w3(32'h3770ff0a),
	.w4(32'h37d71a51),
	.w5(32'h391fe006),
	.w6(32'h380f9c0b),
	.w7(32'h388d6961),
	.w8(32'h3918f336),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c02cb89),
	.w1(32'h3c1daa86),
	.w2(32'h3c0fa956),
	.w3(32'h3c660151),
	.w4(32'h3c421fa9),
	.w5(32'h3bd5f00c),
	.w6(32'h3c8dcdc6),
	.w7(32'h3c36e0da),
	.w8(32'h3c0a5b99),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1a0137),
	.w1(32'hb930991a),
	.w2(32'hb9184aba),
	.w3(32'h3a9ff033),
	.w4(32'h392e5f18),
	.w5(32'hb84f1ba5),
	.w6(32'h3a6e9784),
	.w7(32'h399894d2),
	.w8(32'h39c65f0c),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a598a66),
	.w1(32'hbb3eabf7),
	.w2(32'h3c4aadb8),
	.w3(32'h3c16cc6d),
	.w4(32'hba8060e6),
	.w5(32'h3bbe878b),
	.w6(32'h3c8ecfae),
	.w7(32'h3beda1ea),
	.w8(32'h3be0d3e1),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36b20d1b),
	.w1(32'h374953d1),
	.w2(32'h37d3e055),
	.w3(32'h3726db1a),
	.w4(32'h37467d77),
	.w5(32'h377e86f4),
	.w6(32'h370ff986),
	.w7(32'h3790b4f5),
	.w8(32'h3723b86a),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h369e5ecf),
	.w1(32'h38b3556a),
	.w2(32'h3872d887),
	.w3(32'h381e3bf2),
	.w4(32'h38dc1c5c),
	.w5(32'h3880e1ba),
	.w6(32'h387d2d48),
	.w7(32'h38b9a067),
	.w8(32'h373be76e),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af44213),
	.w1(32'h3b2e935f),
	.w2(32'hbb914033),
	.w3(32'hb81fcf6d),
	.w4(32'h3ab09151),
	.w5(32'hbb6f9ddd),
	.w6(32'hbaed7a3d),
	.w7(32'hb9c14c82),
	.w8(32'hbba1c225),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb34bc1f),
	.w1(32'hba8b4356),
	.w2(32'h39ef6c9a),
	.w3(32'hba97c7c6),
	.w4(32'hbb1a82d0),
	.w5(32'hbadea982),
	.w6(32'h3b04613a),
	.w7(32'hba4659df),
	.w8(32'hba9b8caa),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1824c2),
	.w1(32'h3ac3a5ca),
	.w2(32'hbab58347),
	.w3(32'h3a60710f),
	.w4(32'h392e6eb4),
	.w5(32'hbb1dac1d),
	.w6(32'h3ae393bc),
	.w7(32'h39cfd4f8),
	.w8(32'hbb0d9b25),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b82805e),
	.w1(32'h3c1df35e),
	.w2(32'hba0b36e9),
	.w3(32'hbb00f10e),
	.w4(32'h3b25a0c7),
	.w5(32'hbb801b84),
	.w6(32'hbb1d26f5),
	.w7(32'h38a54ce0),
	.w8(32'hbbfce928),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcce8bf9),
	.w1(32'h3d0edd88),
	.w2(32'h3c21856a),
	.w3(32'hbcbf7ce5),
	.w4(32'h3c8ca89d),
	.w5(32'hbc1d8ab6),
	.w6(32'hbcb3a0d7),
	.w7(32'h3c019a02),
	.w8(32'hbcb5504c),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1c5a43),
	.w1(32'hbc13c6f9),
	.w2(32'h3c0773c8),
	.w3(32'h3bbaa77e),
	.w4(32'hbb4db143),
	.w5(32'h3c0c3607),
	.w6(32'h3cd602b4),
	.w7(32'h3c82c42f),
	.w8(32'h3c242d55),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb84cafd),
	.w1(32'hbc5031d8),
	.w2(32'h3c3f3d16),
	.w3(32'h3c4c05ea),
	.w4(32'hbb7c757f),
	.w5(32'h3c3cbdd8),
	.w6(32'h3cd97198),
	.w7(32'h3c650630),
	.w8(32'h3c91b3c5),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadce693),
	.w1(32'h3a4b5243),
	.w2(32'h3aa04c0b),
	.w3(32'h39f14171),
	.w4(32'h3a96eab0),
	.w5(32'h3affcbeb),
	.w6(32'h3b23604e),
	.w7(32'h3b315654),
	.w8(32'h3aa71232),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3810b2e0),
	.w1(32'h387e81f9),
	.w2(32'h380c6ab2),
	.w3(32'h37fcc36d),
	.w4(32'h3790fdd9),
	.w5(32'hb66ec7fd),
	.w6(32'h37c0c64e),
	.w7(32'h37546c2e),
	.w8(32'hb878b829),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f6221d),
	.w1(32'hb8903e1c),
	.w2(32'h3944d199),
	.w3(32'hb889916c),
	.w4(32'hb82a6d44),
	.w5(32'h392b9503),
	.w6(32'hb46f1be2),
	.w7(32'h3892291f),
	.w8(32'h39095320),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389f575c),
	.w1(32'h3a2a0667),
	.w2(32'h3a88bdfc),
	.w3(32'hb9d2e46e),
	.w4(32'h3a425d4d),
	.w5(32'h37ecba6a),
	.w6(32'h395e359d),
	.w7(32'h3a37b327),
	.w8(32'hb91fa0f6),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0baaa6),
	.w1(32'h3bd7af19),
	.w2(32'hbb8bf6fe),
	.w3(32'h3bb38760),
	.w4(32'h3ba4257b),
	.w5(32'hbb8c9d38),
	.w6(32'hbba4616c),
	.w7(32'hbba195f5),
	.w8(32'hbbaa24d2),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc215d36),
	.w1(32'hbb06cf1f),
	.w2(32'h3b13e1c2),
	.w3(32'hbb916a49),
	.w4(32'h3a5291ce),
	.w5(32'h3b360e05),
	.w6(32'h3aea454c),
	.w7(32'h3baff240),
	.w8(32'h3b97cf03),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1c2b08),
	.w1(32'hba94538c),
	.w2(32'hbb53a3c6),
	.w3(32'hbbdb3325),
	.w4(32'hb93ce390),
	.w5(32'hbba9e1d6),
	.w6(32'hbb99b6b5),
	.w7(32'hba2d26df),
	.w8(32'hbba94f4b),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc0e838),
	.w1(32'hbba1a5d1),
	.w2(32'hbb35cfba),
	.w3(32'hbb5a0430),
	.w4(32'hbb486c55),
	.w5(32'hba2c720a),
	.w6(32'h3a45d37e),
	.w7(32'h3aa82b7f),
	.w8(32'h3a612b5e),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8e9665),
	.w1(32'h3cadc50f),
	.w2(32'hbc1dcdcc),
	.w3(32'h3b7ee2e9),
	.w4(32'h3c0f1f56),
	.w5(32'hbc584ad3),
	.w6(32'hbc2817b6),
	.w7(32'hbb077ca0),
	.w8(32'hbca00afd),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38344983),
	.w1(32'hb88fc8cc),
	.w2(32'hb83ac767),
	.w3(32'h37abefb6),
	.w4(32'hb900a4f3),
	.w5(32'hb609cd3a),
	.w6(32'h37be0567),
	.w7(32'hb87bd220),
	.w8(32'hb881b6ac),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a82dd6),
	.w1(32'hb883c7e2),
	.w2(32'hb9b8baa4),
	.w3(32'hb94f3d15),
	.w4(32'hb87a4085),
	.w5(32'hb9ea166e),
	.w6(32'h37e6e7a1),
	.w7(32'h386ceacb),
	.w8(32'hba044250),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37fc8eb5),
	.w1(32'hb97959ba),
	.w2(32'hb932c0a3),
	.w3(32'h378e5fd8),
	.w4(32'hb9897801),
	.w5(32'hb95e5d49),
	.w6(32'hb909a18c),
	.w7(32'hb9b0b9dd),
	.w8(32'hb99b8f84),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb88976a),
	.w1(32'hbbb0f33b),
	.w2(32'hbb5dfdbf),
	.w3(32'hbbd22077),
	.w4(32'h39cfb1be),
	.w5(32'hbb5eaf0d),
	.w6(32'hbb248f3b),
	.w7(32'hbb087b85),
	.w8(32'hbb23c980),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5ad052),
	.w1(32'h3a51fd18),
	.w2(32'hb8dceabe),
	.w3(32'hbb493137),
	.w4(32'hba8dbaac),
	.w5(32'hb9aa4ed0),
	.w6(32'hbb8a5c7d),
	.w7(32'hbaa3d8e3),
	.w8(32'hbab023de),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c566320),
	.w1(32'h3c4d74af),
	.w2(32'hbc8049dd),
	.w3(32'h3b39a37e),
	.w4(32'h3bd64017),
	.w5(32'hbc6ac465),
	.w6(32'hbb7ec407),
	.w7(32'h3b11ced7),
	.w8(32'hbc84c2f6),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e8506a),
	.w1(32'h3aedfc4d),
	.w2(32'h3a5f6171),
	.w3(32'hb8d1d819),
	.w4(32'h394c93e7),
	.w5(32'h3a1cdcf5),
	.w6(32'hbaad74d2),
	.w7(32'hbaa5a9d9),
	.w8(32'h3ab0d8a4),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91dc795),
	.w1(32'hb734cb14),
	.w2(32'hb88494ba),
	.w3(32'h39a3a4cc),
	.w4(32'hb8874dc0),
	.w5(32'hb9b9f2aa),
	.w6(32'h3a56badb),
	.w7(32'h39639435),
	.w8(32'hb9fbba18),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8052c41),
	.w1(32'h35b4788d),
	.w2(32'hb863718d),
	.w3(32'hb85041ca),
	.w4(32'hb71be192),
	.w5(32'hb887d0c6),
	.w6(32'h37a8c386),
	.w7(32'h37b0672e),
	.w8(32'hb8b70dd2),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398344d1),
	.w1(32'h3a0cc6d7),
	.w2(32'h3aafa87b),
	.w3(32'h3aa4e441),
	.w4(32'h3a4f0bf6),
	.w5(32'h3a8fb0d4),
	.w6(32'h3b12a1fa),
	.w7(32'h3a88d0b7),
	.w8(32'h3a8e6198),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8dd39ba),
	.w1(32'h3a27e24a),
	.w2(32'h3a226b47),
	.w3(32'h39926f26),
	.w4(32'h3a5b8a16),
	.w5(32'h3a3fbb7d),
	.w6(32'h3a3011d1),
	.w7(32'h3a870662),
	.w8(32'h3a289d45),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c0c6bf),
	.w1(32'h3a1c39e5),
	.w2(32'hb9e01181),
	.w3(32'hb8f80b5a),
	.w4(32'h3a1c5973),
	.w5(32'hb9bcda75),
	.w6(32'h3955f00d),
	.w7(32'h3a5b3f72),
	.w8(32'hba657372),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b91c4f1),
	.w1(32'h3b48b6d7),
	.w2(32'hbb9a6fde),
	.w3(32'h38b1ede2),
	.w4(32'h3991f8e0),
	.w5(32'hbbc7be93),
	.w6(32'hbb7e9539),
	.w7(32'hbb3334be),
	.w8(32'hbbd4b59f),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaf8d0b),
	.w1(32'hbbcd983e),
	.w2(32'hbb210e3a),
	.w3(32'hbb4a5168),
	.w4(32'hbb20aa98),
	.w5(32'hbb550247),
	.w6(32'hbbf7acf3),
	.w7(32'hbc178506),
	.w8(32'hbb99b0fc),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7877cf2),
	.w1(32'hb7a9c72d),
	.w2(32'h37bb7142),
	.w3(32'h375e0cb0),
	.w4(32'hb6dfdf10),
	.w5(32'h3474ec18),
	.w6(32'h373c826f),
	.w7(32'hb7a529b8),
	.w8(32'hb7d552bb),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7c5253c),
	.w1(32'h353de5bf),
	.w2(32'h380f59ff),
	.w3(32'h3711bc24),
	.w4(32'h3733a738),
	.w5(32'h37e5d261),
	.w6(32'h37fe0ede),
	.w7(32'h37c8e38b),
	.w8(32'h3787db42),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8121db1),
	.w1(32'hb7f53fc0),
	.w2(32'h37a78205),
	.w3(32'hb85c1a07),
	.w4(32'hb8737bcc),
	.w5(32'hb7ddbbbf),
	.w6(32'hb885d9c3),
	.w7(32'hb7f6491a),
	.w8(32'h36093185),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h386517a9),
	.w1(32'h381e6cb9),
	.w2(32'h38ab85a1),
	.w3(32'h380b205a),
	.w4(32'h37944a67),
	.w5(32'h378499bd),
	.w6(32'h3750ca8b),
	.w7(32'hb772803a),
	.w8(32'hb7786d77),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca215aa),
	.w1(32'h3bdc4a30),
	.w2(32'hbcc1a46a),
	.w3(32'h3c401d35),
	.w4(32'h3aadb4b9),
	.w5(32'hbc9ec69d),
	.w6(32'h3b8324d5),
	.w7(32'hbb0d7f16),
	.w8(32'hbcc2d769),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8eee2a8),
	.w1(32'h3bc29cc8),
	.w2(32'hbb4b1f0c),
	.w3(32'hbbe8038e),
	.w4(32'hbb94c314),
	.w5(32'hbc56251a),
	.w6(32'hbc85339b),
	.w7(32'hbc9152b5),
	.w8(32'hbcc2074d),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb552832),
	.w1(32'hbb7e3cf2),
	.w2(32'hbbf266b5),
	.w3(32'hbb8f32fa),
	.w4(32'hbb472abc),
	.w5(32'hbc10fe63),
	.w6(32'hbbfad480),
	.w7(32'hbc11d096),
	.w8(32'hbbdec20e),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc43909b),
	.w1(32'hbc07c88d),
	.w2(32'h3c1043e3),
	.w3(32'hbb286158),
	.w4(32'hbbe51873),
	.w5(32'h3b5c9330),
	.w6(32'h3c88c63d),
	.w7(32'h3b670c50),
	.w8(32'h3b1a0b17),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37351d9c),
	.w1(32'h38fa278f),
	.w2(32'h38262375),
	.w3(32'h37e95ce2),
	.w4(32'h391144ed),
	.w5(32'hb7769720),
	.w6(32'hb803a233),
	.w7(32'hb6943254),
	.w8(32'hb8a49af0),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h373caf95),
	.w1(32'hb7369f7b),
	.w2(32'h38197891),
	.w3(32'h361ba00f),
	.w4(32'hb8802160),
	.w5(32'hb82cac9c),
	.w6(32'hb7a97057),
	.w7(32'hb812cb0a),
	.w8(32'hb8342897),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3899f2bf),
	.w1(32'hb7830ca1),
	.w2(32'hb6fd0ae5),
	.w3(32'hb737bd79),
	.w4(32'h35b94595),
	.w5(32'hb8a7240d),
	.w6(32'hb82d126b),
	.w7(32'hb90aa689),
	.w8(32'hb9411db7),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5b06e3),
	.w1(32'h3b21096e),
	.w2(32'hbaaa0fb8),
	.w3(32'h3a697cb5),
	.w4(32'h3aaf615a),
	.w5(32'hbaf8f4bc),
	.w6(32'hbb1d1264),
	.w7(32'hbaab9d0a),
	.w8(32'hbb69c9a7),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37afe8a0),
	.w1(32'h38874a8e),
	.w2(32'h38368281),
	.w3(32'h37b26ec4),
	.w4(32'h3851d9ad),
	.w5(32'hb717f1db),
	.w6(32'hb7af4f69),
	.w7(32'hb7eb449d),
	.w8(32'hb85fbf75),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc97440),
	.w1(32'h3c339328),
	.w2(32'hbba962d5),
	.w3(32'h3b59c9e4),
	.w4(32'h3b8736e1),
	.w5(32'hbac558e6),
	.w6(32'hba7065f6),
	.w7(32'h3b9e09d9),
	.w8(32'hbb8ec9ea),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd184bf),
	.w1(32'h3c4e3a5d),
	.w2(32'hbb8e963b),
	.w3(32'hb9288c96),
	.w4(32'h3a6caa06),
	.w5(32'hbbd51ef2),
	.w6(32'hbc354e47),
	.w7(32'hbb3c4d0b),
	.w8(32'hbc6421d6),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc18ae74),
	.w1(32'hbb767b89),
	.w2(32'hba1eff2d),
	.w3(32'hbb6725ef),
	.w4(32'hbb92d379),
	.w5(32'hbad0b6f6),
	.w6(32'h3b4621fd),
	.w7(32'h3b04a03b),
	.w8(32'h3a1fbb69),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b31d946),
	.w1(32'h39a13384),
	.w2(32'hbba6b980),
	.w3(32'hba3713a0),
	.w4(32'hbabcd018),
	.w5(32'hbbb1310b),
	.w6(32'hbb55dde5),
	.w7(32'hbb891618),
	.w8(32'hbbb2de34),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdee614),
	.w1(32'h3c374fcc),
	.w2(32'hbbec56b8),
	.w3(32'h3b2c5c25),
	.w4(32'h3bb8f42a),
	.w5(32'hbc0a5594),
	.w6(32'h3b9a5a16),
	.w7(32'h3ba58c2f),
	.w8(32'hbc174d5d),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbada68ed),
	.w1(32'hbb0ada55),
	.w2(32'h39f76cd7),
	.w3(32'h3aed1d56),
	.w4(32'hba0b65c8),
	.w5(32'hb9d2bac6),
	.w6(32'h3b9edd59),
	.w7(32'h3b1dbd3a),
	.w8(32'h3b0c5fad),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9f5997),
	.w1(32'h3c04afa2),
	.w2(32'hbb277f2f),
	.w3(32'h3aa54498),
	.w4(32'h3b73483f),
	.w5(32'hbb2ea203),
	.w6(32'hbb16cc39),
	.w7(32'h3a560927),
	.w8(32'hbb8872b8),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36269cd2),
	.w1(32'hb7347deb),
	.w2(32'h36ed3fd1),
	.w3(32'h3661a169),
	.w4(32'hb789fa2c),
	.w5(32'hb405b80a),
	.w6(32'hb7829c72),
	.w7(32'hb7d3d8a0),
	.w8(32'hb7277bfa),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3797d68d),
	.w1(32'hb7b6727d),
	.w2(32'hb8aae452),
	.w3(32'h37b6aaa5),
	.w4(32'hb809452f),
	.w5(32'hb881b1a7),
	.w6(32'h390112dc),
	.w7(32'h37c92fc9),
	.w8(32'hb8d43a2b),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb883d622),
	.w1(32'hb8be0401),
	.w2(32'hb8ac1005),
	.w3(32'hb78b1118),
	.w4(32'hb83061d6),
	.w5(32'hb88ad89b),
	.w6(32'hb85b4ede),
	.w7(32'hb74f90e9),
	.w8(32'hb8105f59),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4c3ede),
	.w1(32'h3a9fd810),
	.w2(32'h3a7f5fde),
	.w3(32'h3aee3dd8),
	.w4(32'h3ad71d22),
	.w5(32'h3aba0f82),
	.w6(32'h3b112529),
	.w7(32'h3b0d17f5),
	.w8(32'h3a93d160),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfbbb12),
	.w1(32'hbb3d7ed9),
	.w2(32'h3ab7aaee),
	.w3(32'hbb342dc7),
	.w4(32'hbb5855fd),
	.w5(32'h3a8f8c76),
	.w6(32'h3b7cf752),
	.w7(32'h3b61351f),
	.w8(32'h3b50341a),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a28901),
	.w1(32'h3a4c3593),
	.w2(32'h3a688f6a),
	.w3(32'hb8772068),
	.w4(32'h3a207a4d),
	.w5(32'h39bde96d),
	.w6(32'h39ec9bf0),
	.w7(32'h3a5e55b3),
	.w8(32'h39f3958a),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbae67a2),
	.w1(32'hbb53edfd),
	.w2(32'hbacf4aef),
	.w3(32'hbc01b2e4),
	.w4(32'hbbc22f9b),
	.w5(32'hbb969f38),
	.w6(32'hbb6bc546),
	.w7(32'hbb9c334d),
	.w8(32'hbb95b49f),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0fee90),
	.w1(32'h3c28f7bf),
	.w2(32'hbc0ee96a),
	.w3(32'h3b4d22ab),
	.w4(32'h3b5be071),
	.w5(32'hbbe991f7),
	.w6(32'hbb8e9c50),
	.w7(32'h38e0c6cc),
	.w8(32'hbc1ddbff),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb67f956),
	.w1(32'hbb06c827),
	.w2(32'h3c14b770),
	.w3(32'h3bb9118e),
	.w4(32'h3b58f0ed),
	.w5(32'h3c3885c9),
	.w6(32'h3c65eb93),
	.w7(32'h3c59be55),
	.w8(32'h3c67c3ca),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bec9bc0),
	.w1(32'h3c5961a9),
	.w2(32'hbc68e5b4),
	.w3(32'h3af0b313),
	.w4(32'h3c53bcf4),
	.w5(32'hbc724815),
	.w6(32'h3c028130),
	.w7(32'h3acced4a),
	.w8(32'hbc9cc8cd),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbded846),
	.w1(32'h38001dd1),
	.w2(32'h3b924d7f),
	.w3(32'hbacb279c),
	.w4(32'h3b99d9e0),
	.w5(32'h3c06b889),
	.w6(32'h3b632451),
	.w7(32'h3bfd832a),
	.w8(32'h3c15ff5f),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c34163e),
	.w1(32'h39d18419),
	.w2(32'hbc9404a7),
	.w3(32'h3b43f72a),
	.w4(32'hbbafa307),
	.w5(32'hbcad1ac4),
	.w6(32'hbb277699),
	.w7(32'hbc3b2e50),
	.w8(32'hbcb479c1),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37f8914c),
	.w1(32'hba5ade72),
	.w2(32'hbbe3568b),
	.w3(32'h3b7ce8a4),
	.w4(32'hba2b388c),
	.w5(32'hbb913c5c),
	.w6(32'h3bdfc1b3),
	.w7(32'h3a95a0e6),
	.w8(32'hbb5f92fc),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3993a5ff),
	.w1(32'hbb8aecb6),
	.w2(32'h3bdf3d49),
	.w3(32'h3c13a6d8),
	.w4(32'hba1ea22e),
	.w5(32'h3bbcb53f),
	.w6(32'h3c655e08),
	.w7(32'h3bede4a9),
	.w8(32'h3b9d34b6),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392598f1),
	.w1(32'h395c939b),
	.w2(32'h3980aa67),
	.w3(32'h390659bb),
	.w4(32'h38e2f9de),
	.w5(32'h39873da8),
	.w6(32'h39087987),
	.w7(32'h38ebf428),
	.w8(32'h391e5feb),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3a08de),
	.w1(32'h3b8b1875),
	.w2(32'hbc4216c6),
	.w3(32'hbb46e08c),
	.w4(32'h3afcfe9a),
	.w5(32'hbc36c0e6),
	.w6(32'hbbe70c27),
	.w7(32'hbb6f0a64),
	.w8(32'hbc42980f),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0451f7),
	.w1(32'h3c3472e3),
	.w2(32'hbbe09ea2),
	.w3(32'h3ba0f811),
	.w4(32'h3c290618),
	.w5(32'hbb4dd07e),
	.w6(32'h3c808bcd),
	.w7(32'h3c80dc65),
	.w8(32'hbac42b86),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc62a4e8),
	.w1(32'h3ca41413),
	.w2(32'h3c29282a),
	.w3(32'hbc9f9c70),
	.w4(32'h3b7a13df),
	.w5(32'hbbe2b558),
	.w6(32'hbce5df31),
	.w7(32'hbc3d3d52),
	.w8(32'hbc54ef4a),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0b5385),
	.w1(32'h3bc63a90),
	.w2(32'h3c60ee91),
	.w3(32'h37cb8b10),
	.w4(32'h3c01b29b),
	.w5(32'h3c58b333),
	.w6(32'h3c884fe8),
	.w7(32'h3ca3d798),
	.w8(32'h3c3904d1),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc35a626),
	.w1(32'hbaac1868),
	.w2(32'h3a30a14b),
	.w3(32'hbba5324a),
	.w4(32'hbb330f9d),
	.w5(32'hba8083e0),
	.w6(32'h3b11957b),
	.w7(32'hba843a46),
	.w8(32'hbb1429e7),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c28a58a),
	.w1(32'h3cda5a0a),
	.w2(32'hbbea9ae6),
	.w3(32'hbb348529),
	.w4(32'h3c411a33),
	.w5(32'hbbe36dc0),
	.w6(32'hbb8930eb),
	.w7(32'h3b96a92d),
	.w8(32'hbc4111fa),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a00e9e9),
	.w1(32'h386544f8),
	.w2(32'h36807c9b),
	.w3(32'h39ea7856),
	.w4(32'h3907e4d4),
	.w5(32'h3725e4c5),
	.w6(32'h39f756f3),
	.w7(32'h39255890),
	.w8(32'h370f6ee9),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8c96fd),
	.w1(32'h3c63f452),
	.w2(32'h3bdda198),
	.w3(32'hbc40fa28),
	.w4(32'hbc31da41),
	.w5(32'hbbde2e85),
	.w6(32'hbcb2913b),
	.w7(32'hbbdf61c3),
	.w8(32'hbb3d53eb),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a80957d),
	.w1(32'h3bdc2b3a),
	.w2(32'h3c2cafa2),
	.w3(32'hbb1a7c31),
	.w4(32'h3c0f56b3),
	.w5(32'h3bd8958c),
	.w6(32'hbb04b4f9),
	.w7(32'h3c207be7),
	.w8(32'h3b8d5b71),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38980cbf),
	.w1(32'h393a0f7a),
	.w2(32'h398337a8),
	.w3(32'h37ecb537),
	.w4(32'hb7779aee),
	.w5(32'h38ae8d68),
	.w6(32'h39c97973),
	.w7(32'h39fd54de),
	.w8(32'h39cce95a),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba44f529),
	.w1(32'hbb67ccec),
	.w2(32'hbb38f012),
	.w3(32'h39874fca),
	.w4(32'h39a46cbc),
	.w5(32'hbb9271a1),
	.w6(32'h3b67b711),
	.w7(32'hbaaab64e),
	.w8(32'hbb8531cb),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b151bcf),
	.w1(32'h3bbca737),
	.w2(32'hbbb38f02),
	.w3(32'hba30b1a5),
	.w4(32'h3b75c9a1),
	.w5(32'hbbbec016),
	.w6(32'hbbb5b327),
	.w7(32'hbb1ea57f),
	.w8(32'hbc1213df),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb892dcc),
	.w1(32'hb93763f7),
	.w2(32'h3b17b33d),
	.w3(32'hba9e82e4),
	.w4(32'hba97ec0c),
	.w5(32'h3a449393),
	.w6(32'h3b7dfd45),
	.w7(32'h3b2ab46c),
	.w8(32'h3ad8075d),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb135c40),
	.w1(32'hbbc7847b),
	.w2(32'h3b4a5639),
	.w3(32'h3bc27c40),
	.w4(32'h3a3f825a),
	.w5(32'h3bafc384),
	.w6(32'h3c449839),
	.w7(32'h3baf960c),
	.w8(32'h3c0ae97b),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc102db),
	.w1(32'hbb9b0229),
	.w2(32'hbaa60dd3),
	.w3(32'hbb12f14a),
	.w4(32'hbb5573b5),
	.w5(32'hbae21de7),
	.w6(32'h3aefee99),
	.w7(32'hb88adddb),
	.w8(32'hbaadc727),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b32dfd1),
	.w1(32'h3c3dc5f1),
	.w2(32'h3c019200),
	.w3(32'hbbea9737),
	.w4(32'hba1f5c89),
	.w5(32'hbbbbf354),
	.w6(32'hbb8b3fb5),
	.w7(32'hbbc32cf3),
	.w8(32'hbc31815c),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb8b4d4),
	.w1(32'h3ad773d1),
	.w2(32'hbc2d373e),
	.w3(32'hba333d14),
	.w4(32'hbb114c13),
	.w5(32'hbc2facfd),
	.w6(32'hba8a8e6c),
	.w7(32'hbbcecd7a),
	.w8(32'hbc105c7c),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb45a45f),
	.w1(32'h3a1c51ec),
	.w2(32'h3a5e9e22),
	.w3(32'hba8296a6),
	.w4(32'h3a8ed9e5),
	.w5(32'h3a9db84c),
	.w6(32'h39e5aa96),
	.w7(32'h3adef5f3),
	.w8(32'h3a86770e),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6a38d47),
	.w1(32'hb7c77138),
	.w2(32'hb77e29ad),
	.w3(32'h384a33a3),
	.w4(32'hb83e657b),
	.w5(32'hb89241b0),
	.w6(32'h395ff199),
	.w7(32'h388997ab),
	.w8(32'hb828644d),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9008c10),
	.w1(32'hba3ddfe0),
	.w2(32'hba45335b),
	.w3(32'h38f008da),
	.w4(32'hb72859da),
	.w5(32'hbac1f8b0),
	.w6(32'hb94270fb),
	.w7(32'hba60b8f9),
	.w8(32'hbb1d39c7),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h380ade6f),
	.w1(32'hb8bea721),
	.w2(32'hb80aec31),
	.w3(32'h38204aad),
	.w4(32'hb7cb88b7),
	.w5(32'h369ebb8c),
	.w6(32'hb7ce9803),
	.w7(32'hb79f64fe),
	.w8(32'h3801f9e7),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3938df49),
	.w1(32'hb83a27ed),
	.w2(32'h398f5edc),
	.w3(32'h38f78958),
	.w4(32'h3503a889),
	.w5(32'h398d7b31),
	.w6(32'h38f264c3),
	.w7(32'hb81ef8e9),
	.w8(32'h3894e8ca),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba2c56f),
	.w1(32'hbafbb229),
	.w2(32'hba66a139),
	.w3(32'hbb0c3f9d),
	.w4(32'hb9ce5286),
	.w5(32'hba1dc161),
	.w6(32'h3ab8a925),
	.w7(32'h3a277ea9),
	.w8(32'hb97878f8),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba151ae2),
	.w1(32'h39d3cb63),
	.w2(32'h39dec3ca),
	.w3(32'hb9ae7f93),
	.w4(32'h39a4fdd2),
	.w5(32'h3a288a7c),
	.w6(32'hb96e505d),
	.w7(32'h39cbc4ff),
	.w8(32'h3a095fd0),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdf346e),
	.w1(32'h3bfea2a9),
	.w2(32'hbb829db2),
	.w3(32'h37dd8657),
	.w4(32'h3b4ad39e),
	.w5(32'hbb120edc),
	.w6(32'hbaa3101e),
	.w7(32'h3a8d0206),
	.w8(32'hbbbae0fb),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc8bad9),
	.w1(32'hbc3fa5bf),
	.w2(32'h3b13ceb3),
	.w3(32'h3a563c1b),
	.w4(32'hbc221b72),
	.w5(32'hba9e4166),
	.w6(32'h3c250842),
	.w7(32'hbb511f2a),
	.w8(32'hbaa1b5ae),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c7f126),
	.w1(32'hb89063a5),
	.w2(32'hb88c155a),
	.w3(32'hb86b5d81),
	.w4(32'hb8c49010),
	.w5(32'hb882794d),
	.w6(32'hb7d1b69a),
	.w7(32'hb88c093b),
	.w8(32'hb85342ec),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94f36c6),
	.w1(32'hb954d272),
	.w2(32'hb87f34d6),
	.w3(32'hb58307ca),
	.w4(32'hb88caa95),
	.w5(32'h382b7af0),
	.w6(32'hb721bcdb),
	.w7(32'h364cc12e),
	.w8(32'h385402b3),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h379c4ee1),
	.w1(32'h36b755f5),
	.w2(32'hb68b65a5),
	.w3(32'hb711fe44),
	.w4(32'hb6aa4337),
	.w5(32'hb74178dd),
	.w6(32'hb83d6e56),
	.w7(32'hb7f094cb),
	.w8(32'hb7f5c191),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8adf58),
	.w1(32'hbadd5cba),
	.w2(32'hba61ac59),
	.w3(32'hba1bc399),
	.w4(32'hbbb1e2a8),
	.w5(32'hbb25a7fa),
	.w6(32'h3aa228b1),
	.w7(32'h3bd24b53),
	.w8(32'hbaa5ee8f),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2d6811),
	.w1(32'h3cbc4139),
	.w2(32'hbb4cfb1c),
	.w3(32'hbc2cb294),
	.w4(32'hbb1030ab),
	.w5(32'hbca0bafa),
	.w6(32'hbc2acc3a),
	.w7(32'hbc74d681),
	.w8(32'hbcd8bef6),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2b5843),
	.w1(32'hb9b803d2),
	.w2(32'hbcdf7020),
	.w3(32'h3c003387),
	.w4(32'h3c0cffba),
	.w5(32'hbaf711be),
	.w6(32'hbc729d9b),
	.w7(32'hba023346),
	.w8(32'hbca195d5),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc16fd8),
	.w1(32'h3be8acaf),
	.w2(32'h3bba1897),
	.w3(32'hbc05984a),
	.w4(32'h3bc3bf5b),
	.w5(32'h3bb9e9b5),
	.w6(32'h3ba0ae5c),
	.w7(32'hb9ebadb5),
	.w8(32'h39bd2ad9),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0d2445),
	.w1(32'h3baaf67e),
	.w2(32'hbb3ce6d8),
	.w3(32'h399143e4),
	.w4(32'h37d91a4e),
	.w5(32'hbc2dc94c),
	.w6(32'hbadb2dcc),
	.w7(32'hba801c72),
	.w8(32'hbb4a3835),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8c3217),
	.w1(32'hbc8c1505),
	.w2(32'h3bc7cf41),
	.w3(32'hbb8b1dbf),
	.w4(32'h3bf8b3cb),
	.w5(32'h3bfcafbc),
	.w6(32'h3a501036),
	.w7(32'h3b350a3b),
	.w8(32'h3b218074),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbee335c),
	.w1(32'h3befc929),
	.w2(32'h3a4c029f),
	.w3(32'h3c11edef),
	.w4(32'hbbc2107a),
	.w5(32'hbb762313),
	.w6(32'h3b1aca93),
	.w7(32'hbc706a6f),
	.w8(32'hbc5f6131),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c529447),
	.w1(32'hbc330ea6),
	.w2(32'hbaa52594),
	.w3(32'h3c699608),
	.w4(32'hbb7ec508),
	.w5(32'h3c10f362),
	.w6(32'hba2e5d82),
	.w7(32'hbc31fe74),
	.w8(32'hbc1f7232),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5c0afe),
	.w1(32'h3c6d6465),
	.w2(32'hbc82ebf1),
	.w3(32'h3c1d8b3a),
	.w4(32'h3c2a4003),
	.w5(32'hbc081e62),
	.w6(32'hbb812ab4),
	.w7(32'hbb65b25c),
	.w8(32'hbc78af71),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba481ee3),
	.w1(32'hb9f4a134),
	.w2(32'h3b96e100),
	.w3(32'h3aa117bf),
	.w4(32'hbba61865),
	.w5(32'hbb3eee36),
	.w6(32'h3bde2412),
	.w7(32'h3bad563c),
	.w8(32'h3a77a0e8),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a09d102),
	.w1(32'h3a6ca431),
	.w2(32'hbbf82eaf),
	.w3(32'hbb0ef27d),
	.w4(32'h3af762d2),
	.w5(32'hbba2f7d8),
	.w6(32'hbae99649),
	.w7(32'hbad580bb),
	.w8(32'hbad99cf3),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c632448),
	.w1(32'h3c5c964c),
	.w2(32'hbbbdbc3b),
	.w3(32'h3b687ec1),
	.w4(32'h3c5c3f9e),
	.w5(32'hbb1f3ccf),
	.w6(32'h3a64e95d),
	.w7(32'h391799a0),
	.w8(32'hbbdf1b86),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1390bd),
	.w1(32'hbc8df447),
	.w2(32'hbc8b2a58),
	.w3(32'hbb5dccbd),
	.w4(32'h3a60c4a2),
	.w5(32'h3a52c2e1),
	.w6(32'hbc1be8f4),
	.w7(32'hbc147ae5),
	.w8(32'hbbfced19),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9b1b7e),
	.w1(32'hbba647ac),
	.w2(32'h3b0b2571),
	.w3(32'h38c29c99),
	.w4(32'hbb314d1c),
	.w5(32'hbc372a43),
	.w6(32'hbb7e3d89),
	.w7(32'hbaeb835b),
	.w8(32'hbc685775),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0030a8),
	.w1(32'hba3feb6e),
	.w2(32'hbb5fba95),
	.w3(32'hbb9db100),
	.w4(32'hbb157a2f),
	.w5(32'hbaa02f06),
	.w6(32'h3a17577f),
	.w7(32'h3b8a9347),
	.w8(32'hb689edcb),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8ddf28),
	.w1(32'h3bd3e048),
	.w2(32'h3c4499cc),
	.w3(32'h3c30a7af),
	.w4(32'hbc1c4e81),
	.w5(32'hbcaa6951),
	.w6(32'h3d155bb4),
	.w7(32'h3d1ce0f8),
	.w8(32'h3c501029),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1e3add),
	.w1(32'hbc8a1f56),
	.w2(32'h3c88ce0d),
	.w3(32'hbca719df),
	.w4(32'hbbe7eb18),
	.w5(32'hbcae7b81),
	.w6(32'hbc270ddf),
	.w7(32'hbc85c747),
	.w8(32'hbb0b9270),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc910162),
	.w1(32'h3b02449f),
	.w2(32'h3bc7d074),
	.w3(32'hbc27c094),
	.w4(32'hb909731b),
	.w5(32'h3b1a34d1),
	.w6(32'hbb100ab4),
	.w7(32'hbb9c5526),
	.w8(32'h3a84f7ca),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b58fd4c),
	.w1(32'h3a8013ae),
	.w2(32'hba2e7698),
	.w3(32'h3ae14ef7),
	.w4(32'hbb8d4f4b),
	.w5(32'hbad6a91f),
	.w6(32'hba19b177),
	.w7(32'hbaa12e94),
	.w8(32'hbb9f181b),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb198afe),
	.w1(32'h3b44cd81),
	.w2(32'hba6f3a4f),
	.w3(32'h3a203bf5),
	.w4(32'h3bb0116c),
	.w5(32'h3bad3e1d),
	.w6(32'h3a9442a9),
	.w7(32'hbba5c732),
	.w8(32'h3af5a97d),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdc858c),
	.w1(32'h3b494831),
	.w2(32'h3b3966b5),
	.w3(32'hba386f24),
	.w4(32'h399695f6),
	.w5(32'h39cf11f5),
	.w6(32'h3b10394d),
	.w7(32'h3b8aac3e),
	.w8(32'h3ad83597),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4069de),
	.w1(32'h3bb74438),
	.w2(32'h3a05c791),
	.w3(32'h3a4ee033),
	.w4(32'h3b8d1cb3),
	.w5(32'h39e9f1a7),
	.w6(32'hbafe4b7e),
	.w7(32'hbabf0062),
	.w8(32'hba017da1),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2010c8),
	.w1(32'h3a00c2e1),
	.w2(32'h3b03c488),
	.w3(32'h3b24b105),
	.w4(32'hbb461194),
	.w5(32'hbb80146f),
	.w6(32'hb98a5683),
	.w7(32'h388f38cd),
	.w8(32'hbaf2b36d),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9245bb),
	.w1(32'h3c4270d0),
	.w2(32'hbcb33482),
	.w3(32'hbb0e7cf4),
	.w4(32'hbc119079),
	.w5(32'hbc88113d),
	.w6(32'hbc269d42),
	.w7(32'h3bbddf45),
	.w8(32'hbcae6086),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8750bf),
	.w1(32'h3b9d54c1),
	.w2(32'h393637bd),
	.w3(32'hbc953f49),
	.w4(32'hbb29231e),
	.w5(32'hbb1ac9a6),
	.w6(32'h3a4eecea),
	.w7(32'hbaca404f),
	.w8(32'hbba0fc09),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c42f675),
	.w1(32'h3c60cf72),
	.w2(32'hbc0eec9a),
	.w3(32'hbaa5a781),
	.w4(32'h3bd6696d),
	.w5(32'hbc1119bc),
	.w6(32'h3b8e7c31),
	.w7(32'h3c007b85),
	.w8(32'hbc09d312),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb9709c),
	.w1(32'hbc5f5bd8),
	.w2(32'h3b4ae732),
	.w3(32'h3c069d31),
	.w4(32'h3af8801a),
	.w5(32'h3b552fc1),
	.w6(32'h3cb6fa88),
	.w7(32'h3c14d207),
	.w8(32'h3c42bce5),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd77c7b),
	.w1(32'h3aba8f13),
	.w2(32'h3b15083f),
	.w3(32'hbafa4506),
	.w4(32'h3bb52db3),
	.w5(32'h3b8c5f31),
	.w6(32'h3b9d12b8),
	.w7(32'hbbb6e96d),
	.w8(32'h3a9a85bc),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c10addd),
	.w1(32'h3a87deda),
	.w2(32'h3b3b355a),
	.w3(32'h3b4bb5d9),
	.w4(32'h3a655f46),
	.w5(32'h3b690e39),
	.w6(32'h3a7da235),
	.w7(32'h39e0bee2),
	.w8(32'h3a9d7a71),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5eb7b7),
	.w1(32'h3b273cce),
	.w2(32'h3bde99ed),
	.w3(32'h3af14cbb),
	.w4(32'h3c00bcf7),
	.w5(32'h3bd6a35b),
	.w6(32'h3bd6ab7b),
	.w7(32'hbb9f3166),
	.w8(32'hbb00243d),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b14286),
	.w1(32'hbba9c88c),
	.w2(32'h3bbb96d5),
	.w3(32'h3b560650),
	.w4(32'hbb876f2c),
	.w5(32'h3bf7d836),
	.w6(32'hbb480258),
	.w7(32'h38114deb),
	.w8(32'h3b97a16f),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b23fe8b),
	.w1(32'hbb323247),
	.w2(32'hba74e865),
	.w3(32'h3b5a7c6e),
	.w4(32'hbb9671e2),
	.w5(32'hbb91ac34),
	.w6(32'h3b3de9e4),
	.w7(32'hb88c12c9),
	.w8(32'h3b2a91d1),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c69dc7),
	.w1(32'h3b465e01),
	.w2(32'hbac1f9f2),
	.w3(32'hbb19bb33),
	.w4(32'h3a7979ff),
	.w5(32'hbab44c76),
	.w6(32'h3ae07638),
	.w7(32'h3af6e5fc),
	.w8(32'hbb0b1c31),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf55c98),
	.w1(32'hbb121dd8),
	.w2(32'hbb352615),
	.w3(32'hbac967d6),
	.w4(32'hbad2fa1c),
	.w5(32'hb9ebc221),
	.w6(32'hbb241968),
	.w7(32'hbb553bed),
	.w8(32'hbae54e0a),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2cf0c5),
	.w1(32'h3a0ec9db),
	.w2(32'hbbc68e5c),
	.w3(32'hba81975c),
	.w4(32'hbb8323ac),
	.w5(32'hbc37fba0),
	.w6(32'hbb78608a),
	.w7(32'h3b530216),
	.w8(32'hbbac1c03),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0f6512),
	.w1(32'h3c028b1a),
	.w2(32'h3b30891a),
	.w3(32'h3bed2c1c),
	.w4(32'h3bd4cb0a),
	.w5(32'h3be54112),
	.w6(32'h3b9e7ddb),
	.w7(32'h3ace3f89),
	.w8(32'h3bcf7aa7),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8a5cc7),
	.w1(32'hbb8a609f),
	.w2(32'h3b0e3f5b),
	.w3(32'h3c09da5e),
	.w4(32'h3b4ffd55),
	.w5(32'h3bbce8aa),
	.w6(32'hbadeaea8),
	.w7(32'hbc8106b9),
	.w8(32'hbb600586),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a760bc6),
	.w1(32'hba5b60f2),
	.w2(32'hba8e4b81),
	.w3(32'h3b59bdd4),
	.w4(32'h38dd31e8),
	.w5(32'h39f8ccbc),
	.w6(32'h39dcbe5d),
	.w7(32'hba0e37f4),
	.w8(32'h3ac551f6),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2bf807),
	.w1(32'h3adfdc76),
	.w2(32'h3a6c1061),
	.w3(32'h3b6f1f4d),
	.w4(32'h3bb87726),
	.w5(32'h3b1ee225),
	.w6(32'hba958ffc),
	.w7(32'hbc3beac9),
	.w8(32'hbc25744c),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7f95b7),
	.w1(32'h3b1cecd7),
	.w2(32'hbac20ea4),
	.w3(32'h3b47c0f3),
	.w4(32'h39785557),
	.w5(32'h3a19c6af),
	.w6(32'h39fce5b9),
	.w7(32'hbb0b05c5),
	.w8(32'hbaca7343),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d687ae),
	.w1(32'hb82fbf5e),
	.w2(32'h3b0192dd),
	.w3(32'h36e2c03c),
	.w4(32'h37f5899f),
	.w5(32'h3a46f1aa),
	.w6(32'hbaf8c926),
	.w7(32'hbb0cad19),
	.w8(32'hb9222314),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8630ff),
	.w1(32'hbab39e16),
	.w2(32'h3b404320),
	.w3(32'h3ac5a4e6),
	.w4(32'h39d26c37),
	.w5(32'h3a16de8b),
	.w6(32'h3b80959d),
	.w7(32'h3af7a2b7),
	.w8(32'h3b276f4d),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9f0c7a),
	.w1(32'h3c5df19f),
	.w2(32'hbb8aa744),
	.w3(32'hb9aa3b0b),
	.w4(32'hb9efcaf2),
	.w5(32'hbc239c98),
	.w6(32'hbbe79427),
	.w7(32'h3ae2859b),
	.w8(32'hbbedfdd1),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb923aec5),
	.w1(32'hbc4e23cf),
	.w2(32'hbc95718a),
	.w3(32'hbb572af5),
	.w4(32'hbbeb8044),
	.w5(32'hbc3c18f8),
	.w6(32'hbae935cd),
	.w7(32'hbb94c22c),
	.w8(32'hbbdd9cf3),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca5c145),
	.w1(32'hba74beb2),
	.w2(32'h3b6e5771),
	.w3(32'hbc4396d5),
	.w4(32'hbb68dc74),
	.w5(32'hba00943c),
	.w6(32'h3aa86dcb),
	.w7(32'h3b407d21),
	.w8(32'h3b59ae4e),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cd587e),
	.w1(32'h39b9e5f1),
	.w2(32'hbb692a3c),
	.w3(32'h3b06def7),
	.w4(32'h3bebc1ce),
	.w5(32'h3bb4f818),
	.w6(32'h3b912585),
	.w7(32'h3b0b16b9),
	.w8(32'h3b479990),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc96910),
	.w1(32'hba0515ea),
	.w2(32'hbc978430),
	.w3(32'h3b5daaa1),
	.w4(32'hbb3d925a),
	.w5(32'hbc6e6d4f),
	.w6(32'h3b797f1f),
	.w7(32'h3cbb880b),
	.w8(32'h3c321881),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2d1d53),
	.w1(32'h3b55d7b9),
	.w2(32'hbca06a5a),
	.w3(32'hbbf85e26),
	.w4(32'hbbaeef1d),
	.w5(32'hbc33c6c2),
	.w6(32'h3bffb25d),
	.w7(32'h3ca5f6bd),
	.w8(32'h3b402252),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0cb58d),
	.w1(32'h3b3dc685),
	.w2(32'h3d09f98c),
	.w3(32'hbb758a73),
	.w4(32'h3a353c32),
	.w5(32'hbc49e96d),
	.w6(32'hbc2a6c26),
	.w7(32'hbc6f3f95),
	.w8(32'hbca556a0),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7c5dd9),
	.w1(32'h3ad0742b),
	.w2(32'hbb28e6c1),
	.w3(32'h3b30d2ac),
	.w4(32'h3a90345a),
	.w5(32'h398f982e),
	.w6(32'hbb6c0727),
	.w7(32'hbb8fc5c4),
	.w8(32'h3a8a5b14),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b64957b),
	.w1(32'hbb292b67),
	.w2(32'hbb999310),
	.w3(32'h3b625a69),
	.w4(32'hba523b0a),
	.w5(32'hb99253b6),
	.w6(32'hbac021cf),
	.w7(32'hbb065e79),
	.w8(32'hbb655505),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a950369),
	.w1(32'h3b8f3881),
	.w2(32'h3afa077d),
	.w3(32'h3b00e1cd),
	.w4(32'hbae86723),
	.w5(32'hbbea68f9),
	.w6(32'h3be1a2fc),
	.w7(32'h3c49320e),
	.w8(32'h3b06cd9f),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4030a3),
	.w1(32'h3bcafcfe),
	.w2(32'h3a4b454c),
	.w3(32'hbb9a0ce1),
	.w4(32'hbbb1430c),
	.w5(32'hbca9313e),
	.w6(32'h3c495156),
	.w7(32'h3ca29619),
	.w8(32'h3bba9c0b),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb34e84d),
	.w1(32'hbafe1302),
	.w2(32'h3c8f5ce2),
	.w3(32'hbc23cb44),
	.w4(32'h39f8a1cd),
	.w5(32'hbbd09966),
	.w6(32'hbbd61109),
	.w7(32'hbc95147e),
	.w8(32'hbb8b2d66),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93238bf),
	.w1(32'hbbb53a24),
	.w2(32'h3b9135cb),
	.w3(32'hbc46cc65),
	.w4(32'hbab144ba),
	.w5(32'h3bae3a13),
	.w6(32'hbb917d51),
	.w7(32'hbc3f0b6c),
	.w8(32'hbbec639e),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab68b1a),
	.w1(32'hbb8a683c),
	.w2(32'h3a836b28),
	.w3(32'h39c0eecd),
	.w4(32'hba24197c),
	.w5(32'h3bca455d),
	.w6(32'hbc0ff7ae),
	.w7(32'hbc5dbf75),
	.w8(32'hbb408e34),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c071288),
	.w1(32'hba27f6af),
	.w2(32'h3bb4d440),
	.w3(32'h3bb03c59),
	.w4(32'h3ba091f6),
	.w5(32'h3c23f347),
	.w6(32'hbb8f8543),
	.w7(32'hbbb6bd29),
	.w8(32'hba26dc0b),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4ae9da),
	.w1(32'hbb515dcd),
	.w2(32'hbb79d6d8),
	.w3(32'h3b105417),
	.w4(32'hbbeadc0c),
	.w5(32'hbc04d184),
	.w6(32'h3bc230a2),
	.w7(32'hbad7476c),
	.w8(32'hbabdaf27),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa62aa0),
	.w1(32'h3c612794),
	.w2(32'hbb99807f),
	.w3(32'hbc0283d4),
	.w4(32'h3b5570bb),
	.w5(32'hbc9a6cdc),
	.w6(32'h3cb213a3),
	.w7(32'h3ce699e8),
	.w8(32'h3b8d02c3),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc635287),
	.w1(32'h3c3cec7a),
	.w2(32'h3becf091),
	.w3(32'hbcae2958),
	.w4(32'hbc0b1df2),
	.w5(32'hbc676a3f),
	.w6(32'hbb964e33),
	.w7(32'h3c63e89e),
	.w8(32'hbc67a73e),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf40f20),
	.w1(32'h3b86814f),
	.w2(32'h3b86c145),
	.w3(32'hbc60b544),
	.w4(32'h3b6d6326),
	.w5(32'h3b79be61),
	.w6(32'h3b70ee03),
	.w7(32'hb9b65bc5),
	.w8(32'h3b23b10e),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3bebee),
	.w1(32'h3c1e2724),
	.w2(32'hbc7647c5),
	.w3(32'hba2acc4d),
	.w4(32'h3b2cc2f5),
	.w5(32'hbca92a71),
	.w6(32'hbc2bc400),
	.w7(32'hbbb88f7a),
	.w8(32'hbcadc34a),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8ff515),
	.w1(32'hbc023c2d),
	.w2(32'h3ba9a03c),
	.w3(32'h3c265123),
	.w4(32'hbb8dcd5c),
	.w5(32'h3970016a),
	.w6(32'h3cae312a),
	.w7(32'h3c433d3c),
	.w8(32'h3b6be672),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a425793),
	.w1(32'h3b02b240),
	.w2(32'hbc7be5ea),
	.w3(32'hbabddada),
	.w4(32'hbac7f12d),
	.w5(32'hbbe9723b),
	.w6(32'h3b5ffc8d),
	.w7(32'h3c64bdeb),
	.w8(32'hba492f9a),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbff7368),
	.w1(32'hbaaa6531),
	.w2(32'hbb92ab15),
	.w3(32'hbbf84e06),
	.w4(32'hbb76af20),
	.w5(32'hbb824753),
	.w6(32'hbad101f2),
	.w7(32'h3aa2db63),
	.w8(32'hbb344efc),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8be52d),
	.w1(32'hbac23d25),
	.w2(32'hbb338229),
	.w3(32'h3a86ca7d),
	.w4(32'h3b586085),
	.w5(32'h3b94b22d),
	.w6(32'hb972af9d),
	.w7(32'hbb7941ec),
	.w8(32'h389e3faf),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b21e34c),
	.w1(32'h3b73a78e),
	.w2(32'h3b6aa74a),
	.w3(32'h3b48d305),
	.w4(32'h3bad3585),
	.w5(32'h3bfec490),
	.w6(32'h3a47bb5c),
	.w7(32'h3b1cecad),
	.w8(32'h3ace50c9),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af929b8),
	.w1(32'h3bfdcf2f),
	.w2(32'hbbe21673),
	.w3(32'h3b877298),
	.w4(32'hbb1845d4),
	.w5(32'hbc6707ec),
	.w6(32'h3b267f02),
	.w7(32'h3c860d32),
	.w8(32'hbcb660ff),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc220442),
	.w1(32'hbb072c0f),
	.w2(32'hbc243cdd),
	.w3(32'hbc0035d6),
	.w4(32'hbacbe1df),
	.w5(32'hbbec2e00),
	.w6(32'hbbc12b4a),
	.w7(32'hbb9289a9),
	.w8(32'hbb8683c8),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6b0610),
	.w1(32'hbab08513),
	.w2(32'hba6a9e5f),
	.w3(32'hbc2d9009),
	.w4(32'hbc1ca5b4),
	.w5(32'hbbfcdfda),
	.w6(32'hbb9f3393),
	.w7(32'hbbda65be),
	.w8(32'hbb1c1d4c),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb02de01),
	.w1(32'hbb3cf3f5),
	.w2(32'h3bc1ded5),
	.w3(32'hbbdb2b69),
	.w4(32'hbb4967be),
	.w5(32'hb98a129f),
	.w6(32'hba9047af),
	.w7(32'hbb00d669),
	.w8(32'hb9b20261),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a14b125),
	.w1(32'h3ca3b7a6),
	.w2(32'hbc555430),
	.w3(32'hbb8688cc),
	.w4(32'hbb916db5),
	.w5(32'hbd0f2ace),
	.w6(32'h3c873633),
	.w7(32'h3d0935d6),
	.w8(32'hbbb91d5b),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc13bc6c),
	.w1(32'h3af38c20),
	.w2(32'h3b84adbc),
	.w3(32'hbc7b3990),
	.w4(32'h3b669765),
	.w5(32'h3b92d108),
	.w6(32'hbba936b8),
	.w7(32'hbbf38148),
	.w8(32'hba863a10),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97dddf6),
	.w1(32'h3a674c06),
	.w2(32'h3955c1d5),
	.w3(32'hba6c3a55),
	.w4(32'hba92695f),
	.w5(32'hbb0bb86e),
	.w6(32'h3a4c2cff),
	.w7(32'hba10bea9),
	.w8(32'hbace2585),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b922fdc),
	.w1(32'hbb0310a3),
	.w2(32'hba7113b1),
	.w3(32'h3a4418d0),
	.w4(32'hbbe16439),
	.w5(32'hbb47482d),
	.w6(32'hbbba81bb),
	.w7(32'hbb7ea637),
	.w8(32'hbbb78e23),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bc0a99),
	.w1(32'hbaa94d02),
	.w2(32'hbb1a6b8b),
	.w3(32'h3ab7d360),
	.w4(32'h396f6b72),
	.w5(32'h3ad6e682),
	.w6(32'hbb084ede),
	.w7(32'hbb460d92),
	.w8(32'h399fa04f),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb55e278),
	.w1(32'h3b76f4a3),
	.w2(32'h3b05faa0),
	.w3(32'hba811a97),
	.w4(32'h3b59beae),
	.w5(32'hbaf06a58),
	.w6(32'hbb6c4faf),
	.w7(32'hbb932c59),
	.w8(32'hb947e1d0),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe9f51b),
	.w1(32'hbd10b9a7),
	.w2(32'hb9a98bbc),
	.w3(32'hba5474ee),
	.w4(32'hbcae8732),
	.w5(32'hbce1aa5a),
	.w6(32'h3b0f2a80),
	.w7(32'hbc39f81c),
	.w8(32'hbc1f7b7d),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd04db36),
	.w1(32'h39f18f93),
	.w2(32'hbaa32e2f),
	.w3(32'hbc9f4f67),
	.w4(32'hbb33dff8),
	.w5(32'hbb6de584),
	.w6(32'h3b920d95),
	.w7(32'h3c508c82),
	.w8(32'h3b4cff7f),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3d884f),
	.w1(32'h3a9e4c5b),
	.w2(32'hbb9ac30c),
	.w3(32'hbadb02b6),
	.w4(32'h395430cb),
	.w5(32'hbbf33ff2),
	.w6(32'h3a52f6bc),
	.w7(32'h3b3f1925),
	.w8(32'h3bc456e8),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb80d11),
	.w1(32'hbbaf8c08),
	.w2(32'h3c6244f0),
	.w3(32'hbbffe529),
	.w4(32'h3b1c7a79),
	.w5(32'h3c747c06),
	.w6(32'hbb343fed),
	.w7(32'hbbb9d2f6),
	.w8(32'h3a380b79),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7973eb),
	.w1(32'h3b2b7acb),
	.w2(32'hbb179576),
	.w3(32'h398ec565),
	.w4(32'hba88cbe3),
	.w5(32'hbbf0a24e),
	.w6(32'hba5039b0),
	.w7(32'h3a923a4a),
	.w8(32'hbc0f5ddb),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeeae12),
	.w1(32'h3ba87b0f),
	.w2(32'hba877254),
	.w3(32'h39953d60),
	.w4(32'hba8d8a99),
	.w5(32'hbb8d1139),
	.w6(32'hbb0e017d),
	.w7(32'hbaa6a1f6),
	.w8(32'hbac7b79b),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1599fe),
	.w1(32'h39915d2a),
	.w2(32'hbb2879b6),
	.w3(32'hbb4cbff2),
	.w4(32'hbbc16686),
	.w5(32'hbbd17035),
	.w6(32'h3b7ff23e),
	.w7(32'hbac014ba),
	.w8(32'h3a38c681),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad9a5a2),
	.w1(32'hbb203a25),
	.w2(32'hbb29133e),
	.w3(32'hbc32c35f),
	.w4(32'hbb230180),
	.w5(32'hbbb1254c),
	.w6(32'h3ad60327),
	.w7(32'hbaf920cb),
	.w8(32'h3b115e30),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc140c33),
	.w1(32'h3c1d5c0a),
	.w2(32'hb94a564c),
	.w3(32'hbbddc8e7),
	.w4(32'h3b51dbdc),
	.w5(32'hbb4dcfb6),
	.w6(32'hbbd12b52),
	.w7(32'hbbd2e4ff),
	.w8(32'hbc32d9fc),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b42c3bb),
	.w1(32'h3ac15fd0),
	.w2(32'hbbfbd10d),
	.w3(32'hbb6a89df),
	.w4(32'h3bb43eed),
	.w5(32'hbb4fca95),
	.w6(32'hbc321488),
	.w7(32'hbc1dc940),
	.w8(32'hbc2c73fd),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc310c50),
	.w1(32'hbafbdbde),
	.w2(32'hbba6f778),
	.w3(32'h3a5b7338),
	.w4(32'hbbe41dc6),
	.w5(32'hbc332bec),
	.w6(32'h3b179490),
	.w7(32'h3b48c317),
	.w8(32'hbada539f),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4a9c6c),
	.w1(32'h3cac871c),
	.w2(32'hbc62134d),
	.w3(32'hbbd8e449),
	.w4(32'h3b81673f),
	.w5(32'hbcf3c473),
	.w6(32'h3c996206),
	.w7(32'h3cb3b7aa),
	.w8(32'hbc1bd048),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ada92bd),
	.w1(32'hb990014d),
	.w2(32'hba63a818),
	.w3(32'hbc040740),
	.w4(32'hba62a7ed),
	.w5(32'hbb28858f),
	.w6(32'h3b06c82f),
	.w7(32'hbb1eb937),
	.w8(32'hbb21337e),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a539e5d),
	.w1(32'hba570b9c),
	.w2(32'h3ad5aecb),
	.w3(32'hbadb9a84),
	.w4(32'h3ad3d8a4),
	.w5(32'h3b8f2945),
	.w6(32'hbc12ac73),
	.w7(32'hbc29e51a),
	.w8(32'hbbf3d256),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb741956),
	.w1(32'h3d36fd21),
	.w2(32'h3c39104c),
	.w3(32'hbbcce5e7),
	.w4(32'h3cc0dd30),
	.w5(32'hbc182454),
	.w6(32'hbc5ac8a6),
	.w7(32'h3c5fe3a4),
	.w8(32'hbc8d1314),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be8a1f0),
	.w1(32'h3c241aa2),
	.w2(32'hbc8408bd),
	.w3(32'hbb721f2c),
	.w4(32'h3b2bee06),
	.w5(32'hbc8c8701),
	.w6(32'hbc0ab2da),
	.w7(32'hbbb6c620),
	.w8(32'hbc8962bc),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b338226),
	.w1(32'h3c048070),
	.w2(32'hbc158b56),
	.w3(32'hbaad6610),
	.w4(32'hbb0a77e1),
	.w5(32'hbc39e752),
	.w6(32'hbbd03148),
	.w7(32'h3ae4865c),
	.w8(32'hbc03e9b1),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0dfeab),
	.w1(32'hba99ffa1),
	.w2(32'h3c511e9d),
	.w3(32'hbbf76427),
	.w4(32'h3b2d827e),
	.w5(32'h3ca2235f),
	.w6(32'h3b0ad63e),
	.w7(32'hbbdab741),
	.w8(32'h38b06b00),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe2b85f),
	.w1(32'hbbfadddf),
	.w2(32'h3b149f60),
	.w3(32'h3a7e7c0f),
	.w4(32'hbc1a6c08),
	.w5(32'hbb9fd8fc),
	.w6(32'h3be0e04a),
	.w7(32'hbb3dd0c2),
	.w8(32'hb8c85068),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9ac938),
	.w1(32'h3ae6ed17),
	.w2(32'hba4d1706),
	.w3(32'hbaff7bd2),
	.w4(32'h39e2178c),
	.w5(32'hbae0fb94),
	.w6(32'h3a7711c8),
	.w7(32'h3a47d96b),
	.w8(32'h3a803cac),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a506f98),
	.w1(32'hbb191eb4),
	.w2(32'hbc324558),
	.w3(32'hba75d419),
	.w4(32'hba962ff9),
	.w5(32'h3c6102e0),
	.w6(32'hbc468d48),
	.w7(32'hbb599ee8),
	.w8(32'hbc0f621d),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9bf2b2),
	.w1(32'h3beb1f5b),
	.w2(32'hbabf9d86),
	.w3(32'h3ad90fef),
	.w4(32'hbb85014d),
	.w5(32'hbbe9edd0),
	.w6(32'h3b417925),
	.w7(32'hbb0d0e1b),
	.w8(32'hbbde1e51),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9eca45),
	.w1(32'hba361018),
	.w2(32'hbb492010),
	.w3(32'hbb32e66d),
	.w4(32'h3bba5d24),
	.w5(32'h3c96f142),
	.w6(32'hbba237cd),
	.w7(32'hbc8c1ca4),
	.w8(32'hbaeccf2f),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2a8f39),
	.w1(32'h3be64326),
	.w2(32'h3a6855e6),
	.w3(32'h3c80fd3b),
	.w4(32'h3b2b3cec),
	.w5(32'hba4a2e15),
	.w6(32'h3b93489f),
	.w7(32'h3aaf5650),
	.w8(32'hbb9dfa6f),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af577c6),
	.w1(32'hba6272f6),
	.w2(32'hbbf1b28b),
	.w3(32'hbc0b73a8),
	.w4(32'h3ae2e757),
	.w5(32'hbbb6f75b),
	.w6(32'hbcb72efa),
	.w7(32'hbcf3b037),
	.w8(32'hbcaa6278),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb495cc),
	.w1(32'h3bf5ee2d),
	.w2(32'hbc18c1f2),
	.w3(32'hbb8e00b2),
	.w4(32'hbaf30b76),
	.w5(32'hbc6fac79),
	.w6(32'h3b90fd28),
	.w7(32'h3c89e0a6),
	.w8(32'hbb5c4224),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3fc8a9),
	.w1(32'hbb828f94),
	.w2(32'hbcdcbf12),
	.w3(32'hbc6b3a0d),
	.w4(32'hbbd0dd4c),
	.w5(32'hbbf37aeb),
	.w6(32'h3a389c55),
	.w7(32'hbbfd87be),
	.w8(32'hbc7a49c1),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba13397),
	.w1(32'h3ca8fab9),
	.w2(32'hbba76206),
	.w3(32'hbc6aed52),
	.w4(32'hb85f9430),
	.w5(32'hbc988c55),
	.w6(32'hbb891b22),
	.w7(32'h3c8c9a57),
	.w8(32'hbc69ba2c),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8f198c),
	.w1(32'h3b9f4cfd),
	.w2(32'hbb36999b),
	.w3(32'hbb31a6cc),
	.w4(32'hbaac33ef),
	.w5(32'hbc19e17a),
	.w6(32'hbb066c78),
	.w7(32'hbb4272cd),
	.w8(32'hbc187f34),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b277026),
	.w1(32'h3aa26706),
	.w2(32'hb9feaac1),
	.w3(32'h3b002c88),
	.w4(32'hba889113),
	.w5(32'hbb1afb14),
	.w6(32'h3b4d6a2a),
	.w7(32'h3bde574d),
	.w8(32'h3a310fea),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd319ad),
	.w1(32'h3c2a2158),
	.w2(32'hba6db12c),
	.w3(32'h3b370cfc),
	.w4(32'h3b8ef144),
	.w5(32'hbb41cf95),
	.w6(32'hbaa3ac97),
	.w7(32'h3b1fffcc),
	.w8(32'hbb4e8554),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b360cf2),
	.w1(32'h3b6b5fb2),
	.w2(32'hb9a40b70),
	.w3(32'h3a5d81a4),
	.w4(32'hba56c281),
	.w5(32'hbb504b96),
	.w6(32'h39e2574f),
	.w7(32'h3ac1f468),
	.w8(32'hb8b8422f),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa14977),
	.w1(32'h3a23c87b),
	.w2(32'hba02ff08),
	.w3(32'hbb43ce3f),
	.w4(32'hba8a79c0),
	.w5(32'hbb1c4be2),
	.w6(32'h398c7c9f),
	.w7(32'hba3a2992),
	.w8(32'hbacf3015),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaee40e1),
	.w1(32'h3ae06ba8),
	.w2(32'hbaf81b29),
	.w3(32'hbb0ac6f9),
	.w4(32'hbb260cbf),
	.w5(32'hbb9fd221),
	.w6(32'h3b8f7d0a),
	.w7(32'h3c1cfcb4),
	.w8(32'h3a654ed1),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb375afb),
	.w1(32'h3b52585d),
	.w2(32'h3b13b524),
	.w3(32'hbb143904),
	.w4(32'hba10e693),
	.w5(32'hbc3122e1),
	.w6(32'h3b88507e),
	.w7(32'h3c4aae9a),
	.w8(32'h3be33d71),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb81eff77),
	.w1(32'hb8f4e00b),
	.w2(32'h3c2c0ce4),
	.w3(32'hbbb0573b),
	.w4(32'h3b6306f3),
	.w5(32'h3b90880a),
	.w6(32'hbad9a233),
	.w7(32'hbb81b90c),
	.w8(32'h3b892b07),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c017d49),
	.w1(32'h3bb8688d),
	.w2(32'hbce027b3),
	.w3(32'h3be59e37),
	.w4(32'h3bbe9c50),
	.w5(32'hbcfaeb8e),
	.w6(32'h3b14fbfb),
	.w7(32'h3bfac49b),
	.w8(32'hbb03bf3b),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9148dc),
	.w1(32'h3ba481cd),
	.w2(32'h3adc081d),
	.w3(32'hbc7000d9),
	.w4(32'h3b050656),
	.w5(32'hbbb7126d),
	.w6(32'hbbe90c52),
	.w7(32'hbc0a7986),
	.w8(32'hbc1d418b),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c30b802),
	.w1(32'h3b58d8f9),
	.w2(32'hbcad4f0f),
	.w3(32'h3bfcfb8d),
	.w4(32'h3b2ef0a7),
	.w5(32'hbc96bcb6),
	.w6(32'h3b18f56e),
	.w7(32'h3b246b97),
	.w8(32'hbc234f17),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfd576a),
	.w1(32'h3b576cf9),
	.w2(32'h3b86e944),
	.w3(32'hbbc6b576),
	.w4(32'hbba6aa0f),
	.w5(32'hbc2cec16),
	.w6(32'h3c272ed1),
	.w7(32'h3ca12441),
	.w8(32'h3bb7489e),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8061dd),
	.w1(32'h3aec0959),
	.w2(32'hbb024b8e),
	.w3(32'hbc09f555),
	.w4(32'hbb310144),
	.w5(32'hbbc0fce8),
	.w6(32'h3b9ebed6),
	.w7(32'h3c430138),
	.w8(32'hb990cd7e),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb547305),
	.w1(32'hb943a103),
	.w2(32'hb9e6eddd),
	.w3(32'hbb08c02d),
	.w4(32'hbab98c2e),
	.w5(32'hb9a8a579),
	.w6(32'h3a101352),
	.w7(32'h3b09a331),
	.w8(32'hbaa4d1b0),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb204725),
	.w1(32'hb8fbbdd6),
	.w2(32'h3a19cf36),
	.w3(32'h39e66ae0),
	.w4(32'h3a03f9c2),
	.w5(32'h3b745f34),
	.w6(32'hb951c3f0),
	.w7(32'hb9ca91b0),
	.w8(32'hbae13fe1),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7538b8),
	.w1(32'hbc7f4b36),
	.w2(32'hbd015bf3),
	.w3(32'hbacd1da0),
	.w4(32'hbcb32a91),
	.w5(32'hbcce4a75),
	.w6(32'hbc97b673),
	.w7(32'hbc08b06f),
	.w8(32'hbc9a82cd),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8021a4),
	.w1(32'h3b725b54),
	.w2(32'h39579526),
	.w3(32'hbc512434),
	.w4(32'hbb408d59),
	.w5(32'hbb3cd0ee),
	.w6(32'h3b85b417),
	.w7(32'h3c4ca6cc),
	.w8(32'h3b25d4ff),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa235d6),
	.w1(32'hbb378461),
	.w2(32'h3bb75f6f),
	.w3(32'h3b1b153b),
	.w4(32'h39e8d684),
	.w5(32'h3bdb13fa),
	.w6(32'hb990c2be),
	.w7(32'h3a8dfeea),
	.w8(32'h3b606617),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd7a185),
	.w1(32'hba885be9),
	.w2(32'h3c081323),
	.w3(32'h3bb346b2),
	.w4(32'h3abc394d),
	.w5(32'h3c044608),
	.w6(32'hb97e4359),
	.w7(32'hbb1fca1e),
	.w8(32'hb9d08fec),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc4775d),
	.w1(32'h3ab6742b),
	.w2(32'h399bf970),
	.w3(32'h3bf4d693),
	.w4(32'hba14e240),
	.w5(32'hba5a9f8c),
	.w6(32'h3ad0556c),
	.w7(32'h3b963234),
	.w8(32'h3a65de64),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cbacd4),
	.w1(32'hbc72fc9d),
	.w2(32'hbd224330),
	.w3(32'hb90361c9),
	.w4(32'hbc33594c),
	.w5(32'hbc8e0b2b),
	.w6(32'hbc648c53),
	.w7(32'h390dc974),
	.w8(32'hbca3232c),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca9e21f),
	.w1(32'hbc01e223),
	.w2(32'h3b7427b0),
	.w3(32'hbc80ff04),
	.w4(32'hbb84edca),
	.w5(32'h3c8cb5f6),
	.w6(32'hbc39d23d),
	.w7(32'hbc8cbb97),
	.w8(32'hbc1f2a9e),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bff0411),
	.w1(32'hbb3b181a),
	.w2(32'hbc848ed3),
	.w3(32'h3c2dbf91),
	.w4(32'h3a4e097e),
	.w5(32'hbc513c63),
	.w6(32'hb9b7c10c),
	.w7(32'hbc0d1f0f),
	.w8(32'hbc4548ce),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7634ad),
	.w1(32'h38224df9),
	.w2(32'hbafe784f),
	.w3(32'h39edd779),
	.w4(32'h3acf9106),
	.w5(32'hb9dece75),
	.w6(32'h3aa6849f),
	.w7(32'hb989f3ec),
	.w8(32'hba3c6105),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc12c0f3),
	.w1(32'h3ac57cd4),
	.w2(32'h3b5a651e),
	.w3(32'hbb98721b),
	.w4(32'h38e1ca05),
	.w5(32'hba31f7d3),
	.w6(32'h3aeadde8),
	.w7(32'hbb901cbd),
	.w8(32'hbbd39332),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule