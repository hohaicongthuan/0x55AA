module layer_10_featuremap_456(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0a9484),
	.w1(32'h3a6739e0),
	.w2(32'h3a11c5f0),
	.w3(32'hbabebc34),
	.w4(32'h3a17162a),
	.w5(32'h3a1ce292),
	.w6(32'h39642ab5),
	.w7(32'hb96933c2),
	.w8(32'hba868192),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5d273c),
	.w1(32'hbaece1f8),
	.w2(32'hbb00b69d),
	.w3(32'h3a8ae341),
	.w4(32'hbb1c1440),
	.w5(32'hbae55a29),
	.w6(32'hba5b4baf),
	.w7(32'hbac68264),
	.w8(32'hba8c3c54),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d4fdd3),
	.w1(32'h3a73406d),
	.w2(32'h3850b555),
	.w3(32'h397ce7c2),
	.w4(32'h3a4761db),
	.w5(32'h399ff8a9),
	.w6(32'h36c9fe46),
	.w7(32'h3819d8e7),
	.w8(32'hba184b8b),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac1fd34),
	.w1(32'hbaa78c9f),
	.w2(32'hbacf1399),
	.w3(32'h38da48ae),
	.w4(32'hbaa6568d),
	.w5(32'hba8af1c9),
	.w6(32'hba266e7f),
	.w7(32'hbad1c178),
	.w8(32'h3a808e3c),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac36a50),
	.w1(32'h3a6d66e6),
	.w2(32'h39024ac1),
	.w3(32'hbaa1e0f1),
	.w4(32'h39e3f769),
	.w5(32'h3878e745),
	.w6(32'h3a151c4c),
	.w7(32'hba88a55b),
	.w8(32'hba143afd),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a056496),
	.w1(32'h3a461fec),
	.w2(32'h3ab99c9a),
	.w3(32'hb9a5c087),
	.w4(32'h3a9bbf1f),
	.w5(32'h3a2be637),
	.w6(32'hbac49de4),
	.w7(32'h3a8d84f8),
	.w8(32'h3918cde8),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1756c6),
	.w1(32'h3a9d2dba),
	.w2(32'h38db7af8),
	.w3(32'h3a4fbb47),
	.w4(32'hbac1f663),
	.w5(32'hba503575),
	.w6(32'h3a8219ce),
	.w7(32'h391aeb44),
	.w8(32'hb9b841c2),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba649077),
	.w1(32'h3a1f3557),
	.w2(32'h3a715ffb),
	.w3(32'hbb0d637f),
	.w4(32'hbb03d3a1),
	.w5(32'hbab00922),
	.w6(32'hba0a2708),
	.w7(32'hb9b928ca),
	.w8(32'hb997bf63),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acc39c0),
	.w1(32'hbabfdfc6),
	.w2(32'hbb184c1a),
	.w3(32'h372e9ce8),
	.w4(32'hbb42a336),
	.w5(32'hbb164d11),
	.w6(32'h3abbea5c),
	.w7(32'hbb818aa4),
	.w8(32'hbade42aa),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2cd494),
	.w1(32'h3aff7e2c),
	.w2(32'h3af510cf),
	.w3(32'hbb0670f9),
	.w4(32'h3a640fa2),
	.w5(32'h3a7e5f6b),
	.w6(32'hbb0be035),
	.w7(32'hba032481),
	.w8(32'hba972e32),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8e4aac),
	.w1(32'hbac572ff),
	.w2(32'hba53fdda),
	.w3(32'h393d2edb),
	.w4(32'hba2bb0d2),
	.w5(32'hba4c3dad),
	.w6(32'hba93a5fd),
	.w7(32'hb998f3f4),
	.w8(32'hba32a135),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac18615),
	.w1(32'hba649a31),
	.w2(32'h3984379a),
	.w3(32'hb9f30bf8),
	.w4(32'h3a2a845e),
	.w5(32'h3931a9f1),
	.w6(32'h39e963d2),
	.w7(32'hb6f4df12),
	.w8(32'hb9c28c08),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a83ffbc),
	.w1(32'hba24781f),
	.w2(32'hb9a245f7),
	.w3(32'h3af4b8af),
	.w4(32'hbac62d75),
	.w5(32'hba8009e1),
	.w6(32'h3950ddd4),
	.w7(32'hbb48f541),
	.w8(32'hbb1309f4),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3981d5c1),
	.w1(32'hbaf79602),
	.w2(32'hbabde0d8),
	.w3(32'h38e9730a),
	.w4(32'hbb1c120a),
	.w5(32'hba44913f),
	.w6(32'hba55cc59),
	.w7(32'hba64f858),
	.w8(32'hba521cd9),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96e5f12),
	.w1(32'hba45a419),
	.w2(32'hba4e648c),
	.w3(32'hba9e67f0),
	.w4(32'hbafebd9b),
	.w5(32'hb9db21bd),
	.w6(32'hbad5a5db),
	.w7(32'hbacac136),
	.w8(32'hba66ee90),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4f2a79),
	.w1(32'hb9bc86b8),
	.w2(32'hb8e38b51),
	.w3(32'hbaf02744),
	.w4(32'hbaadcc65),
	.w5(32'hbaf3fd92),
	.w6(32'hb9c118d7),
	.w7(32'hbaad1a35),
	.w8(32'hbaa5ecd8),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a755b2),
	.w1(32'h39ef5d77),
	.w2(32'h39ed6748),
	.w3(32'hbab30e0e),
	.w4(32'h3aa2564b),
	.w5(32'h3acdebb5),
	.w6(32'hbabf370e),
	.w7(32'h3ac97d08),
	.w8(32'h3b1a8251),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2f21d1),
	.w1(32'h3a123bbd),
	.w2(32'h3a610f86),
	.w3(32'h3a4a97da),
	.w4(32'h3a8e68e2),
	.w5(32'h3a8d9d86),
	.w6(32'h3adda2c1),
	.w7(32'h3a0fa8fd),
	.w8(32'hb8cf02ce),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a64fbee),
	.w1(32'hba2eb707),
	.w2(32'hb840ce88),
	.w3(32'h3a03821b),
	.w4(32'hba6efb15),
	.w5(32'h38b9525b),
	.w6(32'hb9612792),
	.w7(32'hbaf8abc7),
	.w8(32'hba6dae36),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91925ef),
	.w1(32'hba29ff3b),
	.w2(32'hb9493b3a),
	.w3(32'hb9936eec),
	.w4(32'h3ab1792e),
	.w5(32'h3a7c446a),
	.w6(32'hba84a68f),
	.w7(32'h39b4ebaa),
	.w8(32'hba51a87b),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafc952b),
	.w1(32'hbacbddeb),
	.w2(32'hba01165f),
	.w3(32'h39c117e0),
	.w4(32'hba908ec8),
	.w5(32'h39eab9ef),
	.w6(32'h39afd44f),
	.w7(32'hbb1fa738),
	.w8(32'hbb1cb2fe),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b3d823),
	.w1(32'hba8fdfb7),
	.w2(32'hbaa83139),
	.w3(32'hb9edb9fa),
	.w4(32'hbae37969),
	.w5(32'hbb2217f9),
	.w6(32'hbac9d67f),
	.w7(32'hbaf51489),
	.w8(32'hbac180f9),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb940c781),
	.w1(32'h38a6224f),
	.w2(32'h3ad4f782),
	.w3(32'hbac76fd2),
	.w4(32'h3af8b015),
	.w5(32'h3b0af461),
	.w6(32'h39136429),
	.w7(32'h3aa1d6c5),
	.w8(32'hb8f0547f),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abb86e5),
	.w1(32'h39937a54),
	.w2(32'hbae81f4a),
	.w3(32'h3b139924),
	.w4(32'hbaf2d7f8),
	.w5(32'hbb546cd5),
	.w6(32'h3ae979bc),
	.w7(32'hbb0836a1),
	.w8(32'hbb61cf48),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8c91a3),
	.w1(32'hb8870d8a),
	.w2(32'h3a204f96),
	.w3(32'hbb3e2055),
	.w4(32'h3a303612),
	.w5(32'h3a4e0cea),
	.w6(32'hbb6f4271),
	.w7(32'hba8e5389),
	.w8(32'hba6925e7),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a8e8c9),
	.w1(32'hba432a34),
	.w2(32'hbab589b6),
	.w3(32'hba8c38ce),
	.w4(32'h39e6c7a5),
	.w5(32'hba15f508),
	.w6(32'hbb30e14e),
	.w7(32'hba8556aa),
	.w8(32'hbab5ce41),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb984f61d),
	.w1(32'hba9d8ad9),
	.w2(32'hbb22896b),
	.w3(32'hba522f8a),
	.w4(32'hbb22cde3),
	.w5(32'hbac10d01),
	.w6(32'hbaa4c87a),
	.w7(32'hbac729b9),
	.w8(32'hbacf8588),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaadd97c),
	.w1(32'h3a55c6ef),
	.w2(32'h3a9116db),
	.w3(32'hbac84017),
	.w4(32'h3a29b90e),
	.w5(32'h3a430013),
	.w6(32'hba6d53fd),
	.w7(32'hb822aa34),
	.w8(32'hba245215),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a022a00),
	.w1(32'hbabc5056),
	.w2(32'hbb16e7da),
	.w3(32'hba81f5aa),
	.w4(32'h3814e76a),
	.w5(32'h37d3f4ea),
	.w6(32'hbaf6cca9),
	.w7(32'hb6974d47),
	.w8(32'hbab2da52),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb022125),
	.w1(32'hbb095b93),
	.w2(32'hb9fe358b),
	.w3(32'hba403b88),
	.w4(32'hb974a0be),
	.w5(32'h39bf93bb),
	.w6(32'hba894752),
	.w7(32'hba468de0),
	.w8(32'hb9adfeeb),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ec49aa),
	.w1(32'hbb3d17a9),
	.w2(32'hba9429da),
	.w3(32'h3a7ff69f),
	.w4(32'hbb2c6c33),
	.w5(32'hba465ab2),
	.w6(32'h39607cd2),
	.w7(32'h3a7e6a21),
	.w8(32'h39c82ca7),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafbe923),
	.w1(32'hba8eb684),
	.w2(32'hbb3604ab),
	.w3(32'hb9da1ed7),
	.w4(32'hbac6d664),
	.w5(32'hbb1016d3),
	.w6(32'hb98d98fc),
	.w7(32'hbae58d8b),
	.w8(32'hbb31023c),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb00e02a),
	.w1(32'h39d26224),
	.w2(32'h39489e0e),
	.w3(32'hbb2790e6),
	.w4(32'hba01bc9c),
	.w5(32'h3aad231e),
	.w6(32'hbb4deef4),
	.w7(32'h380a0196),
	.w8(32'hb95b6d91),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a52bbb9),
	.w1(32'h3aebccfc),
	.w2(32'h3a3a855f),
	.w3(32'hba2c4765),
	.w4(32'h3a983253),
	.w5(32'h3adcb240),
	.w6(32'hba82da36),
	.w7(32'h3a97af5e),
	.w8(32'h3a871168),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96e3833),
	.w1(32'hba2ba1c4),
	.w2(32'hbab3ee77),
	.w3(32'h38acbae5),
	.w4(32'hbab58288),
	.w5(32'hbb1a9195),
	.w6(32'h3a74b768),
	.w7(32'h3967bfcd),
	.w8(32'hb98e2432),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0c3ef3),
	.w1(32'h3a691845),
	.w2(32'h3a249153),
	.w3(32'hbaf31d8a),
	.w4(32'h3942be0d),
	.w5(32'h39608ad2),
	.w6(32'h39baee30),
	.w7(32'hb84c1314),
	.w8(32'h3a637e0f),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3931a44c),
	.w1(32'h38510b39),
	.w2(32'h39126e04),
	.w3(32'h3a326644),
	.w4(32'hb9e3f471),
	.w5(32'h39fc07dd),
	.w6(32'h39894a8a),
	.w7(32'hb986b9ff),
	.w8(32'h3a91c53e),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb915f4bb),
	.w1(32'hbab4039c),
	.w2(32'hbad41719),
	.w3(32'h3a82a826),
	.w4(32'hbb1718b6),
	.w5(32'hbad4f2d6),
	.w6(32'h3b222510),
	.w7(32'hba6fd43e),
	.w8(32'hbae6cb5a),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac04899),
	.w1(32'hba729332),
	.w2(32'hba1920a7),
	.w3(32'hbae0f4df),
	.w4(32'hba8a3d12),
	.w5(32'hb7e16562),
	.w6(32'hbb35f8cd),
	.w7(32'hb9d3cb02),
	.w8(32'hb9208e57),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a98e3f2),
	.w1(32'hb9d5d64d),
	.w2(32'hb9874a30),
	.w3(32'hb7a0a39d),
	.w4(32'h3a19bc01),
	.w5(32'h3a5a2dd0),
	.w6(32'h38d8689b),
	.w7(32'h3a1bad20),
	.w8(32'h39a0290a),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c64d9f),
	.w1(32'hbaa51997),
	.w2(32'hbb5adeed),
	.w3(32'h3a1f1b40),
	.w4(32'hbb19bca0),
	.w5(32'hbb69a43c),
	.w6(32'hb9f42430),
	.w7(32'hbb070e48),
	.w8(32'hbae547ce),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb183980),
	.w1(32'hb9ff673d),
	.w2(32'hba7e83cc),
	.w3(32'hb796ce02),
	.w4(32'hbad49b42),
	.w5(32'hbad674f3),
	.w6(32'hbb1ad4b0),
	.w7(32'hbabc3ec8),
	.w8(32'hbae499ab),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cebf4d),
	.w1(32'h39892186),
	.w2(32'hbafe99df),
	.w3(32'h39abfa8b),
	.w4(32'h3a22dc01),
	.w5(32'hbab8e3bc),
	.w6(32'hb9b4906d),
	.w7(32'h3a4ca672),
	.w8(32'h3a4f0913),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3a19af),
	.w1(32'h3b0a8638),
	.w2(32'h3af46b1f),
	.w3(32'h39014bee),
	.w4(32'h3ac8a31c),
	.w5(32'h3a8ae69b),
	.w6(32'h39c8ff87),
	.w7(32'h3a74eebb),
	.w8(32'h3aca9fac),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb994027d),
	.w1(32'hba4cb889),
	.w2(32'hba06a2f5),
	.w3(32'h37b8f5c6),
	.w4(32'hba4ce5e8),
	.w5(32'h399b98cf),
	.w6(32'h3a613a96),
	.w7(32'hba611ac3),
	.w8(32'hbaa39d68),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99ecef3),
	.w1(32'hba99af3c),
	.w2(32'hba622d9e),
	.w3(32'hba76dff0),
	.w4(32'hbb1f9420),
	.w5(32'hbb780f58),
	.w6(32'hbafd1748),
	.w7(32'hbb030eac),
	.w8(32'hbb11b918),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeb8a0f),
	.w1(32'hbb2ba505),
	.w2(32'hbb40b2e4),
	.w3(32'hbb4786d7),
	.w4(32'hbb13dd98),
	.w5(32'hbb23f362),
	.w6(32'hbb03204c),
	.w7(32'hb9b448aa),
	.w8(32'hb9161c53),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb036db7),
	.w1(32'h39efb4cc),
	.w2(32'h3a8d03d8),
	.w3(32'hbadb94d3),
	.w4(32'hba980e57),
	.w5(32'h39db6092),
	.w6(32'hb95e5bcf),
	.w7(32'h3916f658),
	.w8(32'h3a493f65),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a76799b),
	.w1(32'hbb08884a),
	.w2(32'hbb0c4246),
	.w3(32'h399f4734),
	.w4(32'hbb0a0520),
	.w5(32'hbb24a775),
	.w6(32'h3a12d52d),
	.w7(32'hbb1992d4),
	.w8(32'hbade1fcb),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf98967),
	.w1(32'h39fe8e7e),
	.w2(32'h39f1269c),
	.w3(32'hbb2fa85c),
	.w4(32'h3ad8fdb9),
	.w5(32'h3982933e),
	.w6(32'hbb24c431),
	.w7(32'h3aa3b011),
	.w8(32'hb9ab13a8),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9060c8),
	.w1(32'hb91d6d6f),
	.w2(32'hbadee1f0),
	.w3(32'h3a1deb5d),
	.w4(32'hba680f5e),
	.w5(32'hbb40c82e),
	.w6(32'hbad39a83),
	.w7(32'h386a259b),
	.w8(32'hbb2a248e),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba629040),
	.w1(32'hba9018f4),
	.w2(32'hbab6e232),
	.w3(32'hbacc3548),
	.w4(32'hbafb662b),
	.w5(32'hbb37d003),
	.w6(32'hbb3c1297),
	.w7(32'hbb035083),
	.w8(32'hbacbcec1),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9da0119),
	.w1(32'hba280f81),
	.w2(32'hba57b9c4),
	.w3(32'hba9e66fb),
	.w4(32'hba83821a),
	.w5(32'hba28da68),
	.w6(32'hbaf024b8),
	.w7(32'hba6660ea),
	.w8(32'hbaa0107d),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f65ee4),
	.w1(32'hbb190fbf),
	.w2(32'hbb1cdcb9),
	.w3(32'hba84aac1),
	.w4(32'hbb2ca6ba),
	.w5(32'hbad1c38a),
	.w6(32'hba63a2a0),
	.w7(32'hbb0a9d8f),
	.w8(32'hbb2fe034),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaee001a),
	.w1(32'hb9d03928),
	.w2(32'h38f327b5),
	.w3(32'hbb0ad608),
	.w4(32'hbab75453),
	.w5(32'hbaad2b80),
	.w6(32'hbb36a47a),
	.w7(32'hb9d9a0ee),
	.w8(32'hb94de162),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba56d23c),
	.w1(32'hbaf1dc7b),
	.w2(32'hba3a1e19),
	.w3(32'hbac923c4),
	.w4(32'hbb18ddce),
	.w5(32'hb9ee4186),
	.w6(32'hbaae8626),
	.w7(32'hba034b77),
	.w8(32'hba589392),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f7ddcf),
	.w1(32'hb8cd07c8),
	.w2(32'hb9883ecf),
	.w3(32'hba719877),
	.w4(32'h3958b309),
	.w5(32'hba0c9868),
	.w6(32'hbadfdce7),
	.w7(32'hb9807255),
	.w8(32'hbb10d7ba),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7ec614),
	.w1(32'hba8c9a69),
	.w2(32'hba69bc29),
	.w3(32'hbad304d4),
	.w4(32'hba82b3db),
	.w5(32'hba8602ea),
	.w6(32'hbb1e111f),
	.w7(32'hbae2e11a),
	.w8(32'h3a162434),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaae0786),
	.w1(32'h3a89181a),
	.w2(32'h39c2b4cb),
	.w3(32'hba887eb3),
	.w4(32'h3a68d254),
	.w5(32'hba88c8da),
	.w6(32'hb9598819),
	.w7(32'h3a50dc17),
	.w8(32'h39dab5d0),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb937283e),
	.w1(32'hbb70d916),
	.w2(32'hbb4f9aa8),
	.w3(32'hb99c61c3),
	.w4(32'hbb2eb754),
	.w5(32'hbb0c2956),
	.w6(32'hb97315b2),
	.w7(32'hba3b41dd),
	.w8(32'hba75b595),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba82e2e3),
	.w1(32'hbb70048b),
	.w2(32'hbb6050ab),
	.w3(32'hbb1a3060),
	.w4(32'hbad1b539),
	.w5(32'hba823e94),
	.w6(32'hb98815d9),
	.w7(32'hb96b017b),
	.w8(32'hbaa9b0bc),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1c4a78),
	.w1(32'hba949e21),
	.w2(32'hbab69569),
	.w3(32'hba8f0ae2),
	.w4(32'hba465c6c),
	.w5(32'hb9b5de6e),
	.w6(32'hb9d2fb31),
	.w7(32'hba64988b),
	.w8(32'hbaaa5a6c),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3a9036),
	.w1(32'hba2e90ee),
	.w2(32'hbb014694),
	.w3(32'hba5e9959),
	.w4(32'hbb0337f0),
	.w5(32'hbb2abb55),
	.w6(32'hbac15143),
	.w7(32'hbb2a6f0f),
	.w8(32'hbb4d002c),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf12adf),
	.w1(32'h39a80162),
	.w2(32'h3a90a796),
	.w3(32'hbb34e53b),
	.w4(32'h3aacbae6),
	.w5(32'h3a33db20),
	.w6(32'hbb894680),
	.w7(32'h3aa1458a),
	.w8(32'h39a0267c),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abb33e3),
	.w1(32'h3b4bc45c),
	.w2(32'h3b4d9e9e),
	.w3(32'h3acaea81),
	.w4(32'h3b8490ce),
	.w5(32'h3b89849b),
	.w6(32'h3a725c62),
	.w7(32'h3b6e8f78),
	.w8(32'h3b6b8616),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7d8614),
	.w1(32'h3a3f390a),
	.w2(32'hba0fbfa9),
	.w3(32'h3b8eb11f),
	.w4(32'h3a70d1f3),
	.w5(32'hb7bebc88),
	.w6(32'h3b6aaae4),
	.w7(32'h3a3d3d84),
	.w8(32'h3896c79c),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a17751c),
	.w1(32'h3aa20ff3),
	.w2(32'h3a63120c),
	.w3(32'h3aef44e6),
	.w4(32'h3b0f211d),
	.w5(32'h3ae88559),
	.w6(32'h3aa58eb3),
	.w7(32'h3ad3dc2a),
	.w8(32'h3a3cf5e7),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa15c13),
	.w1(32'h3acf0257),
	.w2(32'h3b1a76cb),
	.w3(32'h3a6fec77),
	.w4(32'h39fe5443),
	.w5(32'h3a97cd8a),
	.w6(32'h3ad92947),
	.w7(32'h38951182),
	.w8(32'hb93dc61a),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac57c3b),
	.w1(32'hba1999c6),
	.w2(32'hbb4a75d9),
	.w3(32'hba992021),
	.w4(32'hbb68f652),
	.w5(32'hbb85da35),
	.w6(32'hbac5527d),
	.w7(32'hbb2a1e2f),
	.w8(32'hbb14f2b8),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb205ecc),
	.w1(32'h3a07b089),
	.w2(32'hbaa64212),
	.w3(32'hbb19b5ba),
	.w4(32'hba5ecb81),
	.w5(32'h3b340f9c),
	.w6(32'hbb1522c4),
	.w7(32'h3992f63d),
	.w8(32'h3a51a95a),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa1f6bf),
	.w1(32'hbaa6f907),
	.w2(32'hba9a2c2d),
	.w3(32'hbaf3a978),
	.w4(32'hba8238ce),
	.w5(32'hbad6edc1),
	.w6(32'hbb40be9c),
	.w7(32'hbae89e6a),
	.w8(32'hbb3fae5a),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac75764),
	.w1(32'hbab04e58),
	.w2(32'hbaf26ab3),
	.w3(32'hbb434162),
	.w4(32'hbb0d8a49),
	.w5(32'hbb3aba74),
	.w6(32'hbb5577cc),
	.w7(32'hba8a2be5),
	.w8(32'hbb9c3f04),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0997b0),
	.w1(32'hb9b9416c),
	.w2(32'h3b7a8ad1),
	.w3(32'hbb049865),
	.w4(32'hbb064f85),
	.w5(32'h3b192e30),
	.w6(32'hbb92b66f),
	.w7(32'hbada20e3),
	.w8(32'h39208c21),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab5b6ab),
	.w1(32'h38f838b7),
	.w2(32'hb9a7f9b9),
	.w3(32'hba2b9804),
	.w4(32'hbab1c4a7),
	.w5(32'hb93eaa4a),
	.w6(32'h3a3a61fd),
	.w7(32'hbb42d210),
	.w8(32'hbb68b8ad),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb393715),
	.w1(32'hbae2ba8a),
	.w2(32'hbaae3fc4),
	.w3(32'hbad451e5),
	.w4(32'hbb93ae94),
	.w5(32'hbb1de182),
	.w6(32'hbb708389),
	.w7(32'hbba5d86d),
	.w8(32'hbaa855a8),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaca0f74),
	.w1(32'hbaed7fae),
	.w2(32'hbb02d398),
	.w3(32'hbb32efd5),
	.w4(32'hbb599bb4),
	.w5(32'hbb076c33),
	.w6(32'hbaac1a4c),
	.w7(32'hbb288d33),
	.w8(32'hbae29f8e),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7be13a),
	.w1(32'h39224a41),
	.w2(32'h398ea1a8),
	.w3(32'hba8ce897),
	.w4(32'h3ae519b8),
	.w5(32'hbb02b79e),
	.w6(32'hbae9cc71),
	.w7(32'hb7bcb349),
	.w8(32'hbab1670f),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba93a31c),
	.w1(32'hbb515ebb),
	.w2(32'hbab64f77),
	.w3(32'hbb9615d5),
	.w4(32'hbbac289f),
	.w5(32'hba4b6f60),
	.w6(32'hbb4d484a),
	.w7(32'hbac98d73),
	.w8(32'hbba54704),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a98aa91),
	.w1(32'h3acfcf0c),
	.w2(32'h394b5b62),
	.w3(32'h3b36d024),
	.w4(32'h3a4e8b8e),
	.w5(32'hbaca8be3),
	.w6(32'hbb97621c),
	.w7(32'h39aa3879),
	.w8(32'h39a5ac11),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afefc72),
	.w1(32'hba8ecc21),
	.w2(32'hbb13e2a9),
	.w3(32'h3ac0597d),
	.w4(32'hb9213497),
	.w5(32'hba40e97c),
	.w6(32'h3b0946d4),
	.w7(32'h3b1bdb09),
	.w8(32'h3b392da9),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f28735),
	.w1(32'h3c1dd72f),
	.w2(32'h3bde3f7d),
	.w3(32'hb9e72796),
	.w4(32'h3bd268da),
	.w5(32'h3b199379),
	.w6(32'h3a2ed4ab),
	.w7(32'h3bdb8a57),
	.w8(32'h3b013bc0),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b89c31b),
	.w1(32'hb9001bcc),
	.w2(32'h3a134f89),
	.w3(32'h3b8f3f59),
	.w4(32'h39570a3f),
	.w5(32'hba43f333),
	.w6(32'h3b2351fc),
	.w7(32'h3b14a6ad),
	.w8(32'hba8c50d2),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b48f582),
	.w1(32'hba3f696d),
	.w2(32'h39a6a3eb),
	.w3(32'hb8a87e49),
	.w4(32'hba2e2703),
	.w5(32'hbae4f45f),
	.w6(32'hba3a7704),
	.w7(32'hba79e5af),
	.w8(32'hbad8d784),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8ea595),
	.w1(32'hba8d4f42),
	.w2(32'hb98afd06),
	.w3(32'hb98d4147),
	.w4(32'hbb08fc14),
	.w5(32'hba9e4353),
	.w6(32'hb9c4f012),
	.w7(32'hbb5d22f0),
	.w8(32'hbbc83c6b),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3959af6e),
	.w1(32'hbabaa910),
	.w2(32'h39078c4f),
	.w3(32'hba9b9177),
	.w4(32'hba4b03f4),
	.w5(32'hbaaa2cec),
	.w6(32'hbba5808b),
	.w7(32'h3b25e49e),
	.w8(32'hbb1583db),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4f5f48),
	.w1(32'hbb6e714c),
	.w2(32'hba02d9e6),
	.w3(32'hbab33c45),
	.w4(32'hbae14529),
	.w5(32'hb9c8ed8f),
	.w6(32'hbb06cf54),
	.w7(32'hbbbe9744),
	.w8(32'hbbac569b),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6c56ca),
	.w1(32'hba8da58c),
	.w2(32'hbb20811c),
	.w3(32'hbbc3d28b),
	.w4(32'hbb148246),
	.w5(32'h3b983f3e),
	.w6(32'hbbbe9dc2),
	.w7(32'hbb411135),
	.w8(32'hba2480a8),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb52093),
	.w1(32'hba4d28d3),
	.w2(32'hbad7ba28),
	.w3(32'h3933a559),
	.w4(32'hbb57d259),
	.w5(32'h3b5d130a),
	.w6(32'h3b16a4e5),
	.w7(32'hbb8b31cf),
	.w8(32'hbb6fad79),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9283e2),
	.w1(32'hbae8cdea),
	.w2(32'hbaa2acdb),
	.w3(32'hba2781e9),
	.w4(32'hbb1b793b),
	.w5(32'hbad6506a),
	.w6(32'h39e07db1),
	.w7(32'hbb29a006),
	.w8(32'hbb088cbe),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa79016),
	.w1(32'hba7510b6),
	.w2(32'hba201b3e),
	.w3(32'hbad23863),
	.w4(32'h3a8f7c5d),
	.w5(32'h3b33de1b),
	.w6(32'hbb39944e),
	.w7(32'hb9770b80),
	.w8(32'h3a5eda84),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b28da45),
	.w1(32'hb9a08c9c),
	.w2(32'hbad509bf),
	.w3(32'h3b39de2a),
	.w4(32'hbac36f0e),
	.w5(32'hbb7b6f55),
	.w6(32'h3b9a84c7),
	.w7(32'hb9837566),
	.w8(32'hbb84f737),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1cc5ec),
	.w1(32'hbb4f096e),
	.w2(32'hba9b7bd6),
	.w3(32'hba4e4412),
	.w4(32'hbb76f5ef),
	.w5(32'hbb0e2ee9),
	.w6(32'hbb0069c5),
	.w7(32'hbb8a924e),
	.w8(32'hbb60cd14),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d82682),
	.w1(32'h3b188637),
	.w2(32'h3ae7620f),
	.w3(32'hb977086f),
	.w4(32'h3a592734),
	.w5(32'hb9d070b6),
	.w6(32'hba0f9a8e),
	.w7(32'h3b338a33),
	.w8(32'hb851faf2),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba358e8b),
	.w1(32'h3ae042ab),
	.w2(32'h3a9870a7),
	.w3(32'hbaa1266b),
	.w4(32'h3b0efa70),
	.w5(32'hb987d405),
	.w6(32'hbafb592d),
	.w7(32'hbabaa329),
	.w8(32'hbb2c8ae8),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa41687),
	.w1(32'hbb69d3ca),
	.w2(32'hbb1334f2),
	.w3(32'h3a9a143d),
	.w4(32'hbaa87553),
	.w5(32'hbb05d10c),
	.w6(32'hbae82699),
	.w7(32'hbb9396b5),
	.w8(32'hbb8ab2e4),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9411e3f),
	.w1(32'h3a060c7f),
	.w2(32'hbb08ec54),
	.w3(32'hb992d45a),
	.w4(32'h3aba340d),
	.w5(32'hbb04afd2),
	.w6(32'hbaf551ee),
	.w7(32'hba0bd435),
	.w8(32'hbb3a0493),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a6c43),
	.w1(32'hbb5bd453),
	.w2(32'hbb2e6cc2),
	.w3(32'hbb7c4dfc),
	.w4(32'hbb7fcfd9),
	.w5(32'hbb861122),
	.w6(32'hbb84d42b),
	.w7(32'hbb369b06),
	.w8(32'hbadaacb8),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb054088),
	.w1(32'hba6c00c7),
	.w2(32'hbac96839),
	.w3(32'hbb80a95a),
	.w4(32'h3b0f7a68),
	.w5(32'h3b360565),
	.w6(32'hbabc7f28),
	.w7(32'h3a6a810c),
	.w8(32'h3b820ac0),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abea935),
	.w1(32'h3a667963),
	.w2(32'h3a981f0f),
	.w3(32'h39e9af35),
	.w4(32'h3a8926c8),
	.w5(32'hb8831fa1),
	.w6(32'hb94f9e7b),
	.w7(32'h3bd97e9a),
	.w8(32'h3b614608),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be21e3c),
	.w1(32'hbba3fe4a),
	.w2(32'hbbb7d060),
	.w3(32'h3be0902b),
	.w4(32'hbb04c92b),
	.w5(32'hba8c4145),
	.w6(32'h3bd821c1),
	.w7(32'hbb408a94),
	.w8(32'hbadce9ee),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6c6dd4),
	.w1(32'hbb2921ca),
	.w2(32'hbb21f95b),
	.w3(32'hb9c99846),
	.w4(32'hbb5f8195),
	.w5(32'hbb311d26),
	.w6(32'hbac33379),
	.w7(32'hbb9485fd),
	.w8(32'hbb49a0ce),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3f75d0),
	.w1(32'h3a518497),
	.w2(32'h3b1f07cf),
	.w3(32'hbb430eb5),
	.w4(32'hb9735b29),
	.w5(32'hba0c6f9a),
	.w6(32'hbb4825df),
	.w7(32'h3ac54a64),
	.w8(32'h3a6728ab),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5df655),
	.w1(32'hb7977940),
	.w2(32'h3a049f52),
	.w3(32'h3aaa9168),
	.w4(32'hba93b976),
	.w5(32'hb919b45b),
	.w6(32'h397d6029),
	.w7(32'hbacead8c),
	.w8(32'hba818c27),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4f3945),
	.w1(32'hb9dabd16),
	.w2(32'hbafe7a4c),
	.w3(32'hbabbb711),
	.w4(32'hba467d43),
	.w5(32'hb94d0f66),
	.w6(32'hbabb5437),
	.w7(32'h3b33c04d),
	.w8(32'h3a11c0e5),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3addc894),
	.w1(32'hba76e710),
	.w2(32'hb964b1ea),
	.w3(32'hba826384),
	.w4(32'hbaacaccc),
	.w5(32'hbb047561),
	.w6(32'hb96815e6),
	.w7(32'hb7e40c70),
	.w8(32'h3abae287),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabb9628),
	.w1(32'hbac81919),
	.w2(32'hba6b8b86),
	.w3(32'hbace614c),
	.w4(32'h3985c9ed),
	.w5(32'hbad3d571),
	.w6(32'h3a27c105),
	.w7(32'hb9bf5362),
	.w8(32'hbad9108b),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398d39c8),
	.w1(32'hbae78d40),
	.w2(32'hba926387),
	.w3(32'hba5cacc1),
	.w4(32'hbb1f501f),
	.w5(32'hbb725208),
	.w6(32'hba8a48dd),
	.w7(32'hbb9b87a6),
	.w8(32'hbb8b3ab2),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3d5917),
	.w1(32'hba3e2d71),
	.w2(32'hba3bedd4),
	.w3(32'hbaa6e3f4),
	.w4(32'hb9eefab8),
	.w5(32'hb9de9c12),
	.w6(32'hbb539ebc),
	.w7(32'h3a0cd844),
	.w8(32'h39f08502),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb93bce5),
	.w1(32'hb9ca9b36),
	.w2(32'hba8f6ced),
	.w3(32'hba7516ee),
	.w4(32'hbb1a9db6),
	.w5(32'hbb14ad3e),
	.w6(32'hba9bf1c5),
	.w7(32'h3b01e77c),
	.w8(32'hb8e3a008),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3978d929),
	.w1(32'hbb64eeda),
	.w2(32'hba6e6d7f),
	.w3(32'hb9b09f96),
	.w4(32'hbb270535),
	.w5(32'h3a0b5d74),
	.w6(32'hbb2b0a45),
	.w7(32'h3b43f129),
	.w8(32'h3b364f91),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac36326),
	.w1(32'hbb3293a7),
	.w2(32'hbb7028b0),
	.w3(32'h39d8bcc8),
	.w4(32'hbb04adca),
	.w5(32'hba85762d),
	.w6(32'h3aff9770),
	.w7(32'h3b3f5a07),
	.w8(32'h3b89a442),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb83e47d),
	.w1(32'hbae4da68),
	.w2(32'hba8001c2),
	.w3(32'h3adc04c4),
	.w4(32'hbaa290c0),
	.w5(32'hbb5cc58d),
	.w6(32'h3b987d09),
	.w7(32'h3a8862c1),
	.w8(32'hbb365feb),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b69128f),
	.w1(32'hbb13c4a8),
	.w2(32'hb99be64c),
	.w3(32'hb70af5ab),
	.w4(32'hbad67eaa),
	.w5(32'hbaeefba3),
	.w6(32'hbb1fb3f0),
	.w7(32'hbb5be6b9),
	.w8(32'hbb78ea44),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5cc6ca),
	.w1(32'h3abdb0b3),
	.w2(32'h3b0c8197),
	.w3(32'hbb72b7cb),
	.w4(32'hba900c31),
	.w5(32'h3ab27655),
	.w6(32'hbb19894e),
	.w7(32'hbb33102c),
	.w8(32'hba9026a8),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb05eee6),
	.w1(32'h39068ea4),
	.w2(32'h39f5ba0a),
	.w3(32'hbb4283f3),
	.w4(32'h3b3579f7),
	.w5(32'h3bd8d4b0),
	.w6(32'hbb63d5dd),
	.w7(32'h3a3c6dff),
	.w8(32'h3b91caa9),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb79a470),
	.w1(32'h3ace108a),
	.w2(32'h38ac1add),
	.w3(32'hb960ce4b),
	.w4(32'h3adc7a2e),
	.w5(32'hba37c589),
	.w6(32'h3b28567c),
	.w7(32'h3ac8a5b9),
	.w8(32'hbaca588a),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa6ae2b),
	.w1(32'h3aad78ee),
	.w2(32'h3b8e3e1f),
	.w3(32'h3a79ad06),
	.w4(32'hb9137d0a),
	.w5(32'h3b72cea3),
	.w6(32'h3a987228),
	.w7(32'hbaef23e4),
	.w8(32'h3adc7028),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac9e00e),
	.w1(32'h3ae58072),
	.w2(32'h389494cf),
	.w3(32'h3b018dcd),
	.w4(32'h3a7ed7a8),
	.w5(32'hba9651c8),
	.w6(32'h3b4a35d2),
	.w7(32'h3b363032),
	.w8(32'h3a3d99fa),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b82bc52),
	.w1(32'h3a47de7c),
	.w2(32'hb9de3a5b),
	.w3(32'h3b5f85e2),
	.w4(32'hbb51e810),
	.w5(32'h3a10762b),
	.w6(32'h3a37cd48),
	.w7(32'hbb2fc870),
	.w8(32'hbb029789),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba965d52),
	.w1(32'hbaef3edd),
	.w2(32'h3ab1025f),
	.w3(32'h3b00c096),
	.w4(32'hbb1327d2),
	.w5(32'hb9cc3462),
	.w6(32'hbb3a97c1),
	.w7(32'hbb7df5bd),
	.w8(32'hba9cf4f9),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7a3633),
	.w1(32'h3a96b3bd),
	.w2(32'hb9da0cfc),
	.w3(32'h3a40a93b),
	.w4(32'h3ae2f7aa),
	.w5(32'hbb6df831),
	.w6(32'h3a72bd4e),
	.w7(32'h3a8e4b40),
	.w8(32'hba6c06c5),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf5e7c7),
	.w1(32'hba805614),
	.w2(32'hbbcfb07f),
	.w3(32'hbb5f4cc9),
	.w4(32'hbaf49b5b),
	.w5(32'hbb03e027),
	.w6(32'hbae47096),
	.w7(32'hbb298479),
	.w8(32'hba4c8b19),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2afae3),
	.w1(32'hbae36db0),
	.w2(32'hba48e0da),
	.w3(32'hb8492e8f),
	.w4(32'hbb283f2b),
	.w5(32'hbb59a888),
	.w6(32'hbb10a0a7),
	.w7(32'hbb8e2fbf),
	.w8(32'hbb669eea),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9c8585),
	.w1(32'h3af5f68b),
	.w2(32'h3bdc156d),
	.w3(32'hbb44de2a),
	.w4(32'h3b5118a6),
	.w5(32'h3a7f6c09),
	.w6(32'hbaa55708),
	.w7(32'h3a7f4947),
	.w8(32'h3a49615a),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc0fb5d),
	.w1(32'hbb006091),
	.w2(32'h3b33f1d5),
	.w3(32'h3b481d0a),
	.w4(32'hbb531312),
	.w5(32'h39fbb183),
	.w6(32'h39c78693),
	.w7(32'hba346c4e),
	.w8(32'hbacaec5c),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8f8473),
	.w1(32'hba7916c8),
	.w2(32'hbab62eb3),
	.w3(32'h3b3cb218),
	.w4(32'hbb4c3153),
	.w5(32'hbb140ad2),
	.w6(32'hbade0701),
	.w7(32'h38dbf404),
	.w8(32'h3aab5f7e),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeaea5d),
	.w1(32'hbb7413f6),
	.w2(32'hba72de28),
	.w3(32'hbb32f2e7),
	.w4(32'hbb8d5505),
	.w5(32'h3a33fc5b),
	.w6(32'h3a0af350),
	.w7(32'hbb7538f1),
	.w8(32'hbaf11e21),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9e40d4),
	.w1(32'hba4fad3b),
	.w2(32'h37d78010),
	.w3(32'h392ee8bb),
	.w4(32'hba76ed7a),
	.w5(32'hb8b0bf2d),
	.w6(32'hb90ef6f1),
	.w7(32'hbb009c71),
	.w8(32'hbb001d46),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1bc009),
	.w1(32'hb9db7c3c),
	.w2(32'h3a63413d),
	.w3(32'hbaf51880),
	.w4(32'h3942674a),
	.w5(32'h3b237bc6),
	.w6(32'hb99b2736),
	.w7(32'h3ad304ea),
	.w8(32'h3b2f0531),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390d1c79),
	.w1(32'hb9c11de6),
	.w2(32'hbb07603d),
	.w3(32'h3b9b014f),
	.w4(32'hbacd118b),
	.w5(32'hba80bb07),
	.w6(32'h3b7d5fe8),
	.w7(32'hbae34d05),
	.w8(32'hbb16b24c),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb19e268),
	.w1(32'hbb637420),
	.w2(32'hba007cea),
	.w3(32'hbaaa9c1b),
	.w4(32'hbb2b8d09),
	.w5(32'h3b2932b4),
	.w6(32'hbaa5b143),
	.w7(32'hbb3a3205),
	.w8(32'hb9748eb3),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba212a0e),
	.w1(32'hbabd28ab),
	.w2(32'hbab94316),
	.w3(32'h3a4ea449),
	.w4(32'hbba83b7d),
	.w5(32'hbb182ea3),
	.w6(32'h3b040164),
	.w7(32'hbb1267ee),
	.w8(32'h3a58e0d3),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb094a22),
	.w1(32'hb98e1270),
	.w2(32'hba7fc5e8),
	.w3(32'h39f3cd03),
	.w4(32'hbb000fcb),
	.w5(32'hbb6c0405),
	.w6(32'h39600c70),
	.w7(32'hba7b6c2f),
	.w8(32'hbad60d70),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9674b0),
	.w1(32'hba9e9194),
	.w2(32'h3ac76a71),
	.w3(32'hbb16af62),
	.w4(32'h3b0bc3cb),
	.w5(32'h3acafc67),
	.w6(32'hba66c8be),
	.w7(32'h3aba2e15),
	.w8(32'h3b3a6cba),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9bfb96),
	.w1(32'h3b181a6b),
	.w2(32'h3adcde82),
	.w3(32'h3a1398d6),
	.w4(32'hbb532f03),
	.w5(32'h394d1b98),
	.w6(32'hbaad5e5d),
	.w7(32'hbafaaf5c),
	.w8(32'hbb8084d4),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a32934f),
	.w1(32'h3a4927ef),
	.w2(32'h3b3f1d30),
	.w3(32'h3a9ce6a0),
	.w4(32'hb98c2ae1),
	.w5(32'hb9a8053d),
	.w6(32'hbb5aafbd),
	.w7(32'hbb4429ca),
	.w8(32'hbb1736f6),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afd6a38),
	.w1(32'h3a263c8d),
	.w2(32'hba50054e),
	.w3(32'h3b415d54),
	.w4(32'hba3546d7),
	.w5(32'h3a819863),
	.w6(32'hbb2548da),
	.w7(32'hb988ea41),
	.w8(32'hba1f6f54),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb20a660),
	.w1(32'h3a70f06c),
	.w2(32'h3ae74be3),
	.w3(32'hba48ee4c),
	.w4(32'h3828e37f),
	.w5(32'h3a1f791c),
	.w6(32'hbb00c57d),
	.w7(32'h39cb0984),
	.w8(32'hb9c3a6da),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4f4baa),
	.w1(32'hba9c3de7),
	.w2(32'h3a25910a),
	.w3(32'h3af78ef1),
	.w4(32'hbb02157f),
	.w5(32'hbadd17bd),
	.w6(32'hba58fee1),
	.w7(32'hb9a8c85e),
	.w8(32'hba917cf5),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8913f3),
	.w1(32'h3ac55da8),
	.w2(32'h3aef73e1),
	.w3(32'h3997e582),
	.w4(32'h3a8c39d6),
	.w5(32'hba926412),
	.w6(32'h3971e3fd),
	.w7(32'hb92c7db3),
	.w8(32'hbb287dcf),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b578d4d),
	.w1(32'hbb86dd65),
	.w2(32'hbb50d38a),
	.w3(32'hbac9fa29),
	.w4(32'hbadb3982),
	.w5(32'hbbb6ad18),
	.w6(32'hbb0851f5),
	.w7(32'hbb4e4d04),
	.w8(32'hbba38e46),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h384cf71a),
	.w1(32'hbae7ff1f),
	.w2(32'hbabf77cb),
	.w3(32'hbba0fce1),
	.w4(32'hba91b284),
	.w5(32'hb87fd68d),
	.w6(32'hbbb07181),
	.w7(32'h3a0a5876),
	.w8(32'hba2fa643),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb18d378),
	.w1(32'hbadf2748),
	.w2(32'h39a03e78),
	.w3(32'hba698742),
	.w4(32'hba91165d),
	.w5(32'h360b37cb),
	.w6(32'hbaee8a88),
	.w7(32'h3a923037),
	.w8(32'hbaf54880),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a09bf77),
	.w1(32'hba49aa9f),
	.w2(32'hb9beb0e8),
	.w3(32'hb982ae0c),
	.w4(32'h364100cb),
	.w5(32'hbab1f368),
	.w6(32'hbab8d046),
	.w7(32'h39bd008f),
	.w8(32'hbb3c561e),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94afa91),
	.w1(32'h3af3490d),
	.w2(32'h3b38adbf),
	.w3(32'h3960a983),
	.w4(32'hb9a6ac60),
	.w5(32'h3aed7736),
	.w6(32'hbac6b241),
	.w7(32'h3ae44f64),
	.w8(32'h3a834f96),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aae73da),
	.w1(32'h3b77076e),
	.w2(32'h3b2160c3),
	.w3(32'h3b62fb34),
	.w4(32'h3b1293d9),
	.w5(32'h3b60ca91),
	.w6(32'h3b233d00),
	.w7(32'h3afbedef),
	.w8(32'h3b469dff),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a90c0f0),
	.w1(32'hbb135874),
	.w2(32'h39a11624),
	.w3(32'h3afc87c3),
	.w4(32'hbb91e343),
	.w5(32'hbb86607a),
	.w6(32'h3b918bdc),
	.w7(32'hba8961b3),
	.w8(32'hbadbf435),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af2b8c7),
	.w1(32'h3a76abc9),
	.w2(32'hbadd5124),
	.w3(32'h39d8d727),
	.w4(32'hba3ffa24),
	.w5(32'hba3f7d47),
	.w6(32'h3812f1c1),
	.w7(32'h3b83c9c1),
	.w8(32'h3a81aeca),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae22829),
	.w1(32'h3afa8b6a),
	.w2(32'h3b0ccc86),
	.w3(32'hbabdd0e4),
	.w4(32'h3b807c45),
	.w5(32'h3abacc4c),
	.w6(32'h3b18ca98),
	.w7(32'h3a87121e),
	.w8(32'h3a938e70),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b417d09),
	.w1(32'h39f6145d),
	.w2(32'hb9ca2234),
	.w3(32'hbad2252c),
	.w4(32'h3a69d9f9),
	.w5(32'h3b99ae8b),
	.w6(32'hba574848),
	.w7(32'h3a19c2df),
	.w8(32'h3b62354d),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb176ab9),
	.w1(32'hbb7ca491),
	.w2(32'hbaea6731),
	.w3(32'hba617d13),
	.w4(32'hbb1cf301),
	.w5(32'h39e53f23),
	.w6(32'hba490265),
	.w7(32'h389357aa),
	.w8(32'hba0f8bc4),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb49ddae),
	.w1(32'h3ab2eb61),
	.w2(32'hb9852a72),
	.w3(32'h3ade9d74),
	.w4(32'hb9f4d5ca),
	.w5(32'hbb4798e2),
	.w6(32'hba543e74),
	.w7(32'h3aa6d497),
	.w8(32'hba5a91a9),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba14d368),
	.w1(32'hbb1a04e7),
	.w2(32'hbb279550),
	.w3(32'hbb3feac3),
	.w4(32'hbb1b812a),
	.w5(32'hba834aca),
	.w6(32'hbaa517c4),
	.w7(32'hbb1c359b),
	.w8(32'hbb46f05e),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1805b7),
	.w1(32'h3b65deff),
	.w2(32'hbab08b91),
	.w3(32'hbaca0fc7),
	.w4(32'h3b98b794),
	.w5(32'h3b1484e1),
	.w6(32'hbab010dc),
	.w7(32'h3af1980c),
	.w8(32'hba42cdd3),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb37565e),
	.w1(32'hba419065),
	.w2(32'h3addb785),
	.w3(32'hbacd37ef),
	.w4(32'hba494aa5),
	.w5(32'h3a7de6a2),
	.w6(32'hbb889d0e),
	.w7(32'h3b59aeb3),
	.w8(32'h3bb9283b),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b440b71),
	.w1(32'h3aa05e33),
	.w2(32'hba55f6de),
	.w3(32'h3b6b9200),
	.w4(32'hb9f7ea7a),
	.w5(32'hb9c8b312),
	.w6(32'h3bb766fb),
	.w7(32'h3a867986),
	.w8(32'hba106220),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2e1c8b),
	.w1(32'hb9bc337d),
	.w2(32'hb8c5ac90),
	.w3(32'hbaadd9f6),
	.w4(32'hbb3abe58),
	.w5(32'hbb0454eb),
	.w6(32'hbaa28aee),
	.w7(32'hbb406cc8),
	.w8(32'hbb2520d4),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba54feb7),
	.w1(32'hbb5e4b2c),
	.w2(32'hbb180cd9),
	.w3(32'hbb2c8d67),
	.w4(32'hbb13bea0),
	.w5(32'hbb809b29),
	.w6(32'h399ed480),
	.w7(32'h394842e4),
	.w8(32'hbb06f8dd),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a76cfc0),
	.w1(32'hb99cf2ca),
	.w2(32'hb9845f86),
	.w3(32'hbb4b60cf),
	.w4(32'hbb6a2043),
	.w5(32'hbb00e4ff),
	.w6(32'hbb8afa36),
	.w7(32'hbb72cbf5),
	.w8(32'hbb5c094e),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b02b5af),
	.w1(32'hbb5b7eba),
	.w2(32'h39b0aaaa),
	.w3(32'hbaa52e9b),
	.w4(32'hbb272a9e),
	.w5(32'h3a8e8293),
	.w6(32'hbaa36698),
	.w7(32'hbb8d39ee),
	.w8(32'hbae150c0),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a858db1),
	.w1(32'h3ae4fe70),
	.w2(32'hba2c4e02),
	.w3(32'h3b1e3149),
	.w4(32'h3b219e3f),
	.w5(32'h3a1cff25),
	.w6(32'h3ad30aff),
	.w7(32'h3a43bf02),
	.w8(32'hbaf9635e),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1c58d0),
	.w1(32'h3ae9ff8c),
	.w2(32'hbafb9611),
	.w3(32'hbb4a39ff),
	.w4(32'h3a9652bb),
	.w5(32'hba8b65b2),
	.w6(32'hbb838712),
	.w7(32'h3b07852c),
	.w8(32'hbb447392),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaba5c69),
	.w1(32'h3b1f2144),
	.w2(32'h3abc13ad),
	.w3(32'h3a3c1452),
	.w4(32'h3b5c38ea),
	.w5(32'h3949dc4e),
	.w6(32'hbb4095cf),
	.w7(32'h3bb4f9dd),
	.w8(32'h3a759511),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b836478),
	.w1(32'h3ae6df26),
	.w2(32'h3a2b8c06),
	.w3(32'h3b4f3827),
	.w4(32'h3a839975),
	.w5(32'h3ae86b97),
	.w6(32'hba7e983d),
	.w7(32'h3a83f528),
	.w8(32'h3ae3dac2),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba66c9b0),
	.w1(32'hbae426be),
	.w2(32'hba5b6a75),
	.w3(32'h3a9d04f7),
	.w4(32'hbb054025),
	.w5(32'hbafcf447),
	.w6(32'h3a3ba7df),
	.w7(32'hba86f815),
	.w8(32'hbb1693d2),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3f79aa),
	.w1(32'hbb0c9a99),
	.w2(32'hba860610),
	.w3(32'hbac16c29),
	.w4(32'hbb547450),
	.w5(32'hbb39bed0),
	.w6(32'hbb15e142),
	.w7(32'hbb826f4e),
	.w8(32'hbbaba990),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392354ab),
	.w1(32'h3b67e1de),
	.w2(32'h3b6ec10f),
	.w3(32'hba603890),
	.w4(32'h3b9a6c36),
	.w5(32'h3b93ccaa),
	.w6(32'hbb7defc6),
	.w7(32'h3b5c2f82),
	.w8(32'h3b4ea338),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba457a30),
	.w1(32'h3a6971d3),
	.w2(32'h3a593b7a),
	.w3(32'h3b3080ff),
	.w4(32'hbb505bf9),
	.w5(32'h3b03aae7),
	.w6(32'h3b86ff55),
	.w7(32'hbb3749be),
	.w8(32'hba91d4ab),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa35c39),
	.w1(32'hbb61d624),
	.w2(32'hbb30cb93),
	.w3(32'h3b8593eb),
	.w4(32'hbb079be4),
	.w5(32'hbb8dbbc1),
	.w6(32'h3ae04841),
	.w7(32'hbb43aee1),
	.w8(32'hbb3e79e3),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7a38f2),
	.w1(32'hba800298),
	.w2(32'h3ade40f6),
	.w3(32'hbbcbe3cf),
	.w4(32'hba9ee38e),
	.w5(32'hbaa5d01b),
	.w6(32'hbba9ddd1),
	.w7(32'hbaa1ee18),
	.w8(32'h3a0f7082),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0ca86e),
	.w1(32'h39d85ec3),
	.w2(32'h3a815202),
	.w3(32'h3932c05b),
	.w4(32'hb8cf4341),
	.w5(32'h3a9b4081),
	.w6(32'h3a5523e6),
	.w7(32'h39bb387f),
	.w8(32'h3b248fcc),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae1f16c),
	.w1(32'h3b09745b),
	.w2(32'h3b900c3c),
	.w3(32'h3b5ba140),
	.w4(32'h3b3cb287),
	.w5(32'h3bc016ff),
	.w6(32'h3b95665f),
	.w7(32'h3b1ab883),
	.w8(32'h3b827610),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b74a6fc),
	.w1(32'h3b1173e2),
	.w2(32'h3b3fa2ed),
	.w3(32'h3c0f3fa7),
	.w4(32'hba2eada8),
	.w5(32'hb93c9858),
	.w6(32'h3c0a73fb),
	.w7(32'hb8115a2b),
	.w8(32'h373e4136),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cd7024),
	.w1(32'hbaa91634),
	.w2(32'hbb848809),
	.w3(32'hbaef690c),
	.w4(32'hbb0f0164),
	.w5(32'hbb3e7098),
	.w6(32'hbaf47899),
	.w7(32'hbab83a6c),
	.w8(32'hbbc5cf7f),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb673f04),
	.w1(32'hbb6a748a),
	.w2(32'hbb011e27),
	.w3(32'hbb794b72),
	.w4(32'hbaea5a2f),
	.w5(32'h3ae4c462),
	.w6(32'hbb780ab6),
	.w7(32'hbae73ba1),
	.w8(32'h3a3a3a3b),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb661adf),
	.w1(32'hbb211e16),
	.w2(32'hbb246745),
	.w3(32'hba32979d),
	.w4(32'hbb13e372),
	.w5(32'hbb2c793d),
	.w6(32'h3a9e925d),
	.w7(32'hba99603e),
	.w8(32'hbb3c55da),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2d6ba5),
	.w1(32'h3979b627),
	.w2(32'hbae845c4),
	.w3(32'hbae9303d),
	.w4(32'hba10049f),
	.w5(32'hbad67cae),
	.w6(32'hbaaf0222),
	.w7(32'h3b2cad75),
	.w8(32'h3a084576),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2d6b7c),
	.w1(32'hbb81dbf6),
	.w2(32'h3a18df52),
	.w3(32'hbabfe02d),
	.w4(32'hbb253d15),
	.w5(32'hbb104832),
	.w6(32'hba880667),
	.w7(32'hbbc35b95),
	.w8(32'hbb4c01eb),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a871d0d),
	.w1(32'hbace46ee),
	.w2(32'hbb305b91),
	.w3(32'h3af136df),
	.w4(32'hb72131e1),
	.w5(32'hbb142264),
	.w6(32'h3a3dc006),
	.w7(32'h3ad5f2bf),
	.w8(32'h3aab9e0b),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaacbe88),
	.w1(32'hbaf43f8b),
	.w2(32'hbb2dc6e8),
	.w3(32'hbb5b969d),
	.w4(32'hbb49d969),
	.w5(32'h39eaaf0b),
	.w6(32'hbae54b3d),
	.w7(32'hba927fe1),
	.w8(32'h3ad08b99),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6997ad),
	.w1(32'h3b39b561),
	.w2(32'h3af61314),
	.w3(32'hbb2fdbda),
	.w4(32'h3aec2169),
	.w5(32'h3b13ff38),
	.w6(32'hba62b295),
	.w7(32'h39f97cb2),
	.w8(32'hbaa638c7),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38baa819),
	.w1(32'h3b1f8369),
	.w2(32'h39b3da57),
	.w3(32'hb90c2422),
	.w4(32'h3b06f3cb),
	.w5(32'h3af94ac1),
	.w6(32'hbb02c96c),
	.w7(32'h3a8331ad),
	.w8(32'hba925f5f),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0c8d89),
	.w1(32'hba9e9738),
	.w2(32'h3b30baab),
	.w3(32'hbb2b6ba5),
	.w4(32'hbaf0aa71),
	.w5(32'h3b78e1fa),
	.w6(32'hbb4d50c1),
	.w7(32'h3b1fafb4),
	.w8(32'h3af0ae8f),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb25c00a),
	.w1(32'h3afd1a19),
	.w2(32'hba030b92),
	.w3(32'h3b8e894a),
	.w4(32'h3aba2076),
	.w5(32'h3b4f582b),
	.w6(32'h3ba41900),
	.w7(32'h3b0300af),
	.w8(32'h3a83e66d),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaf5254),
	.w1(32'hba825d7d),
	.w2(32'h3ae78894),
	.w3(32'h37e75e54),
	.w4(32'h37941616),
	.w5(32'hbada5a01),
	.w6(32'h3a7b5061),
	.w7(32'h3ac430ea),
	.w8(32'h3b731641),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf70140),
	.w1(32'hbafb201a),
	.w2(32'hbb324a43),
	.w3(32'h3bc22305),
	.w4(32'h3a82e54f),
	.w5(32'hba2d48ca),
	.w6(32'h3bd55c75),
	.w7(32'hb9327016),
	.w8(32'h3b394275),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3add84a7),
	.w1(32'hbbad9d13),
	.w2(32'hbb254fa8),
	.w3(32'hbaadff5f),
	.w4(32'hbba4fa54),
	.w5(32'hba108939),
	.w6(32'hb8e5446c),
	.w7(32'hbb85603a),
	.w8(32'h38d847bb),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb12f015),
	.w1(32'hb9c2d822),
	.w2(32'hba5281bd),
	.w3(32'hba75f345),
	.w4(32'hbb6348a4),
	.w5(32'h3aa55367),
	.w6(32'h3a5d3239),
	.w7(32'hbbae40f4),
	.w8(32'hbb90a85a),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb510a40),
	.w1(32'h3ab27bd7),
	.w2(32'h3abe1db4),
	.w3(32'h3abfa19a),
	.w4(32'hb9b3d835),
	.w5(32'h3b04f02f),
	.w6(32'h3b1df43f),
	.w7(32'h3b87abbc),
	.w8(32'h3bb34585),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba590f06),
	.w1(32'h3909671c),
	.w2(32'h3b7ac2b1),
	.w3(32'h3b8a029e),
	.w4(32'h3a694adc),
	.w5(32'h393eebe4),
	.w6(32'h3c356a2d),
	.w7(32'h3b1dc696),
	.w8(32'h3882649a),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95a2e50),
	.w1(32'hbb5b1708),
	.w2(32'hb88f1e5d),
	.w3(32'h3b2723f5),
	.w4(32'hbb26d6ba),
	.w5(32'h3b03e60b),
	.w6(32'h3b0ef770),
	.w7(32'hbb3d7693),
	.w8(32'h3ac9d765),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a65a73),
	.w1(32'h3a4ac7c5),
	.w2(32'h3a328448),
	.w3(32'h3b1f9fbe),
	.w4(32'hb9df887f),
	.w5(32'hbb3d5a56),
	.w6(32'h3b98e523),
	.w7(32'h3a479f84),
	.w8(32'h3a9596ca),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b763219),
	.w1(32'h3b7a9255),
	.w2(32'h3b2cfaf8),
	.w3(32'h390bdf12),
	.w4(32'h3b1c39d6),
	.w5(32'h3a9f2010),
	.w6(32'h3b00197a),
	.w7(32'h3b3710fa),
	.w8(32'h3b14b6b7),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8fc3a0),
	.w1(32'h3bb58fc2),
	.w2(32'h3b0ae3e1),
	.w3(32'h3ba06447),
	.w4(32'h3bbd6d92),
	.w5(32'h3a761cdf),
	.w6(32'h3b995516),
	.w7(32'h3b8260a8),
	.w8(32'hb918fac4),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae8f0dd),
	.w1(32'h398eca94),
	.w2(32'hb9955d3e),
	.w3(32'hbace3738),
	.w4(32'h3ad4910c),
	.w5(32'h3b07eec6),
	.w6(32'hbac014f4),
	.w7(32'h39b47b73),
	.w8(32'h39db9ac4),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3938259d),
	.w1(32'hbb2a562e),
	.w2(32'hbb3f5639),
	.w3(32'h3ab9ec23),
	.w4(32'hbb0eb6e1),
	.w5(32'hbbe3111b),
	.w6(32'h3aab24de),
	.w7(32'h3a0aca62),
	.w8(32'hbb4ba611),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb75faee9),
	.w1(32'hbb155f01),
	.w2(32'hbaeb73c0),
	.w3(32'hbb24e8ed),
	.w4(32'hbb121928),
	.w5(32'hba0d57bd),
	.w6(32'hbaf34d58),
	.w7(32'hbb0478b1),
	.w8(32'hbafa2104),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb97b28a),
	.w1(32'h3b5958e4),
	.w2(32'h3b733e4b),
	.w3(32'hbba2b01b),
	.w4(32'hba808258),
	.w5(32'hbb17d7f2),
	.w6(32'hbb92071d),
	.w7(32'hb9a65218),
	.w8(32'hbb452367),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1fd238),
	.w1(32'hba2de21a),
	.w2(32'h3b54f5d6),
	.w3(32'h3b9c4b5c),
	.w4(32'h3c2e46d1),
	.w5(32'h3c4e5ceb),
	.w6(32'h3c3c9386),
	.w7(32'h3bcc7332),
	.w8(32'h3a8e9622),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba027482),
	.w1(32'h3b37fcd3),
	.w2(32'h3a20c6b3),
	.w3(32'h3ab598f3),
	.w4(32'hbc3b4627),
	.w5(32'hbc7ad071),
	.w6(32'h3aa3c039),
	.w7(32'hbbac9024),
	.w8(32'h3a0c11ec),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb515d84),
	.w1(32'hbb97eae7),
	.w2(32'hbb9d0214),
	.w3(32'hbbdf3b42),
	.w4(32'h3b6418f5),
	.w5(32'h3a5082ad),
	.w6(32'h3b8b7463),
	.w7(32'h3bd5b90d),
	.w8(32'hbb28c1aa),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8dfefe),
	.w1(32'h3b667846),
	.w2(32'hbabec1d8),
	.w3(32'h3b605a28),
	.w4(32'h396f7430),
	.w5(32'hbad709d9),
	.w6(32'hbad6c103),
	.w7(32'h3a5b869c),
	.w8(32'hb9c8e9f5),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadee061),
	.w1(32'hbbd7a4c5),
	.w2(32'h3abf7084),
	.w3(32'h38bc4028),
	.w4(32'hbba9e5ae),
	.w5(32'h3b2b24a8),
	.w6(32'hbb8ed897),
	.w7(32'h3a8a320a),
	.w8(32'hbadaf8ec),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad37f9f),
	.w1(32'h3acf14c1),
	.w2(32'hbb088245),
	.w3(32'hbbf189d7),
	.w4(32'h399f6462),
	.w5(32'hbbcab21b),
	.w6(32'hbc1928c3),
	.w7(32'h3b06ad57),
	.w8(32'h3acfb843),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7a939d8),
	.w1(32'h3c7b767c),
	.w2(32'h3c1971c7),
	.w3(32'hba5a4279),
	.w4(32'h3b1cd1a7),
	.w5(32'h3ca72066),
	.w6(32'h37a04a65),
	.w7(32'hbb7459d1),
	.w8(32'h3c9f8c59),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3c9961),
	.w1(32'hbc163f4a),
	.w2(32'hbc10625a),
	.w3(32'h3c4527b3),
	.w4(32'hbc114f37),
	.w5(32'hbc4b9029),
	.w6(32'h3c1aa7e3),
	.w7(32'hbb262fa2),
	.w8(32'hbbed1c0f),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b01dc94),
	.w1(32'h3a23f301),
	.w2(32'h3b467155),
	.w3(32'hbbeb6b71),
	.w4(32'h3a7663f0),
	.w5(32'h3ab38f3a),
	.w6(32'hbc06f6a1),
	.w7(32'h3bc969df),
	.w8(32'h3a856c94),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0e497a),
	.w1(32'h3c370fb6),
	.w2(32'h3c92090a),
	.w3(32'h3b0b3983),
	.w4(32'h3a71d416),
	.w5(32'h3d254643),
	.w6(32'h3b88f020),
	.w7(32'hbace47b5),
	.w8(32'hbba39c2b),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1f35d4),
	.w1(32'h3bda178a),
	.w2(32'h3b80ac68),
	.w3(32'h3bf2467e),
	.w4(32'h3bd14338),
	.w5(32'hba4d1f6c),
	.w6(32'h3c2b3c33),
	.w7(32'h3b80d864),
	.w8(32'h3bdbe1c8),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9537a3),
	.w1(32'h3b826f1d),
	.w2(32'h3b840bca),
	.w3(32'h3bba7908),
	.w4(32'h3ae2cd4f),
	.w5(32'hbb29552a),
	.w6(32'h3b8c610a),
	.w7(32'h3a8afc9a),
	.w8(32'hb9d49b91),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8424b8),
	.w1(32'hbb8fe837),
	.w2(32'hbbf73638),
	.w3(32'h3b611cc1),
	.w4(32'h3b6d0e79),
	.w5(32'hbac3675d),
	.w6(32'hbadd3935),
	.w7(32'h3ae0d30c),
	.w8(32'hbb9fe91b),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb95bf3),
	.w1(32'hbb2ea90c),
	.w2(32'h3bd24d2f),
	.w3(32'h3b3125b6),
	.w4(32'h3c598562),
	.w5(32'h3c53c2bd),
	.w6(32'hba61a701),
	.w7(32'h3c3e9a4e),
	.w8(32'hbb9786c2),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bffdb17),
	.w1(32'h399f1817),
	.w2(32'h3b262411),
	.w3(32'h3c19abd6),
	.w4(32'h3ab58db7),
	.w5(32'hbb02643e),
	.w6(32'hbb054907),
	.w7(32'h3bb5b8f2),
	.w8(32'h3bc82b7e),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf3ea21),
	.w1(32'hba4da20a),
	.w2(32'hbbb13c65),
	.w3(32'hbaecb10f),
	.w4(32'h3c1f7b44),
	.w5(32'hbc03f6df),
	.w6(32'hbb57999f),
	.w7(32'hbb114610),
	.w8(32'hbbb2e094),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba72d216),
	.w1(32'hbbdb0be4),
	.w2(32'hba9a8c1d),
	.w3(32'h3a244a2d),
	.w4(32'h3a62a578),
	.w5(32'h3cd1f175),
	.w6(32'h3a46788c),
	.w7(32'h3baa16b7),
	.w8(32'h3ae8b154),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h375be3fe),
	.w1(32'hbbbc4d82),
	.w2(32'hbbf836df),
	.w3(32'h3c00580f),
	.w4(32'hbb562d8b),
	.w5(32'h3c4a0816),
	.w6(32'hbb0caee2),
	.w7(32'h3b6a2c55),
	.w8(32'h3b30fca7),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbce926e),
	.w1(32'h3c10ee95),
	.w2(32'h3bfdd83f),
	.w3(32'hbb1197b3),
	.w4(32'h3bf1d524),
	.w5(32'h3c832d78),
	.w6(32'hbb9c3952),
	.w7(32'h3a6c66cf),
	.w8(32'h3c078848),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3e8463),
	.w1(32'hbb6adde0),
	.w2(32'hb8461342),
	.w3(32'h3b99d7a8),
	.w4(32'hbafec190),
	.w5(32'hba9fa432),
	.w6(32'h3a2159fa),
	.w7(32'h3b886b6d),
	.w8(32'hbabf778f),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa95ecf),
	.w1(32'hba6d4536),
	.w2(32'hbbdb9396),
	.w3(32'hbb66799b),
	.w4(32'h3b235f39),
	.w5(32'h3addbb8b),
	.w6(32'hbb8f66eb),
	.w7(32'h3a9d8ec1),
	.w8(32'h3b90c647),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb044bdc),
	.w1(32'hba5b240a),
	.w2(32'hbba155ff),
	.w3(32'hbba43cc8),
	.w4(32'h3c2dcc61),
	.w5(32'h3c6c3bc2),
	.w6(32'hbb6f45ec),
	.w7(32'h3b9295dd),
	.w8(32'hba8a2cd5),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbea7bce),
	.w1(32'h3a060f5d),
	.w2(32'hb9c280b8),
	.w3(32'h3c190d6e),
	.w4(32'h3a8b472d),
	.w5(32'hb904a774),
	.w6(32'h3664ec5d),
	.w7(32'hba5d23e8),
	.w8(32'hbb06045c),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaad599),
	.w1(32'hbb86bb70),
	.w2(32'hbc0bddaf),
	.w3(32'h3b2f30b3),
	.w4(32'h3a6257d2),
	.w5(32'hbbdc5aca),
	.w6(32'h3b918e0a),
	.w7(32'hba36643a),
	.w8(32'hbac252b3),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc06d260),
	.w1(32'h3ae6e084),
	.w2(32'hb98ec6ba),
	.w3(32'hbb6cfd58),
	.w4(32'h3c33b6c6),
	.w5(32'h3cc20a91),
	.w6(32'h3acec4ed),
	.w7(32'hb9324c1e),
	.w8(32'hb92c033d),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb310ed6),
	.w1(32'h3a8c00c7),
	.w2(32'hbba249da),
	.w3(32'hbb1e49c7),
	.w4(32'hbc07e4a4),
	.w5(32'hba52f1d2),
	.w6(32'hbb467ca4),
	.w7(32'hbbe95ff2),
	.w8(32'hba7a7501),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc641b5),
	.w1(32'h3b7298db),
	.w2(32'hbb088231),
	.w3(32'hbbe901c2),
	.w4(32'h3b69831b),
	.w5(32'hbb3a1f07),
	.w6(32'hbb3cce3f),
	.w7(32'hb9c93cbe),
	.w8(32'h3a9dd658),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a578723),
	.w1(32'h3b0a414d),
	.w2(32'h3b098b71),
	.w3(32'h3b90cd94),
	.w4(32'h3b01f835),
	.w5(32'h3b59d644),
	.w6(32'h3b39d160),
	.w7(32'hbae10bb8),
	.w8(32'hbabff284),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3c1108),
	.w1(32'hb93d4422),
	.w2(32'h3b01bc4d),
	.w3(32'h3ba19014),
	.w4(32'h3b4fd485),
	.w5(32'h3be1cd07),
	.w6(32'hbb02c586),
	.w7(32'h3ab8a9c0),
	.w8(32'h3b479782),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9948d4),
	.w1(32'hbc340e84),
	.w2(32'hbbd06827),
	.w3(32'h3aea9ba7),
	.w4(32'hbbaac727),
	.w5(32'hbb8c08f7),
	.w6(32'hbba2a959),
	.w7(32'h3abc5709),
	.w8(32'h393427cc),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb52a351),
	.w1(32'h3b540733),
	.w2(32'hb9973884),
	.w3(32'hbbfcda0f),
	.w4(32'h3c4de730),
	.w5(32'h3c5b3021),
	.w6(32'hbbfd5b18),
	.w7(32'h3aed7c54),
	.w8(32'h3c095e61),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8459a93),
	.w1(32'hbb8a13c4),
	.w2(32'hbbdd7872),
	.w3(32'h3b09a74c),
	.w4(32'hbae1c29b),
	.w5(32'hb8b96c98),
	.w6(32'h3b7c239d),
	.w7(32'hb9ecbecd),
	.w8(32'hb913e07a),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3d2659),
	.w1(32'hbb26fa5c),
	.w2(32'hbb8b68f8),
	.w3(32'hbbb26118),
	.w4(32'h3a5e7d62),
	.w5(32'hbc24ffbd),
	.w6(32'hbb95bbd1),
	.w7(32'h3bbc4226),
	.w8(32'hbb859f5f),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa4e67e),
	.w1(32'hbc1cc5f5),
	.w2(32'hbbd98a8f),
	.w3(32'hbb8fd63a),
	.w4(32'hbc2d3779),
	.w5(32'hbc18eaf4),
	.w6(32'hbb4eb233),
	.w7(32'hbb62faaf),
	.w8(32'hbb548b29),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac2cb4c),
	.w1(32'hbaf8343c),
	.w2(32'hbbcc598b),
	.w3(32'hbb2d76d4),
	.w4(32'h3bc26a46),
	.w5(32'h3bd069eb),
	.w6(32'hbb75d8ae),
	.w7(32'hbb0df116),
	.w8(32'hbb923493),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc4484d),
	.w1(32'h39882184),
	.w2(32'hbb70b9c5),
	.w3(32'h3b9f8424),
	.w4(32'h3be4b9b1),
	.w5(32'hb8b704f2),
	.w6(32'h3bb72f6c),
	.w7(32'hba925e0b),
	.w8(32'h3a9efb92),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0d774c),
	.w1(32'h3b14f928),
	.w2(32'h3b5cb6c5),
	.w3(32'hbb93abd3),
	.w4(32'h3bb2c1e9),
	.w5(32'hb9b7f09e),
	.w6(32'h3b30eafe),
	.w7(32'h3a9dd98f),
	.w8(32'hbb6d62c9),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaae3f77),
	.w1(32'h3a8f99b5),
	.w2(32'hba5c8c03),
	.w3(32'hba11f59a),
	.w4(32'hbb2818f0),
	.w5(32'h38b104db),
	.w6(32'hbb98f980),
	.w7(32'h3b37c0f9),
	.w8(32'hbadd6397),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b92bc1d),
	.w1(32'hbb1ee6c4),
	.w2(32'hbb2c4d3e),
	.w3(32'hbb17bb1c),
	.w4(32'h399e20f5),
	.w5(32'hb98e74c8),
	.w6(32'hbb99badd),
	.w7(32'hbb4b629d),
	.w8(32'hbb918320),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9b242b),
	.w1(32'hbb9eb736),
	.w2(32'hbc40b5d0),
	.w3(32'hbb978fe3),
	.w4(32'h3b081e7d),
	.w5(32'h3ca0ef80),
	.w6(32'hba980bcb),
	.w7(32'hbb184a60),
	.w8(32'hbb8384b0),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb7fff0),
	.w1(32'hbb6c7b4d),
	.w2(32'h3ae93960),
	.w3(32'hbb0f3b65),
	.w4(32'h3bc0e84e),
	.w5(32'h3a22f022),
	.w6(32'h3a3a501c),
	.w7(32'hbab09b80),
	.w8(32'h3a827267),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad9322f),
	.w1(32'hbb137d7d),
	.w2(32'hbb76cf15),
	.w3(32'h3b21be76),
	.w4(32'hbb059fa7),
	.w5(32'hbc01c14f),
	.w6(32'h3a5d6fa1),
	.w7(32'hbc1106b7),
	.w8(32'hbb90a669),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1bff12),
	.w1(32'hbada0592),
	.w2(32'hbc00c288),
	.w3(32'hbbec90eb),
	.w4(32'hbb225917),
	.w5(32'hbaa27f07),
	.w6(32'hbbf97274),
	.w7(32'h3b076bbd),
	.w8(32'h3b3417dc),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f0182),
	.w1(32'h3ba2fa3a),
	.w2(32'h3b04d5c1),
	.w3(32'h3a661452),
	.w4(32'hba593150),
	.w5(32'hbc1f5d0e),
	.w6(32'hba741970),
	.w7(32'hbb10e231),
	.w8(32'hbc080951),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcdadc8),
	.w1(32'hbc04d140),
	.w2(32'hbc1d3987),
	.w3(32'h3ad82441),
	.w4(32'hbbbe69bb),
	.w5(32'hbbd436a5),
	.w6(32'hbaf92e06),
	.w7(32'hbab80bc0),
	.w8(32'hbbcf4bd3),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc25c971),
	.w1(32'hbbcf2606),
	.w2(32'hbb0803e5),
	.w3(32'hbab7f99c),
	.w4(32'h3a91e22a),
	.w5(32'hbb366f00),
	.w6(32'hbb18c4ef),
	.w7(32'h3c142142),
	.w8(32'hbb8f499e),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4edc5b),
	.w1(32'hba485625),
	.w2(32'hbc27e0b3),
	.w3(32'hbba08d89),
	.w4(32'h39c0cc6f),
	.w5(32'hb93ea051),
	.w6(32'hbb051f94),
	.w7(32'h3aad5ff7),
	.w8(32'h3a1566b0),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf62854),
	.w1(32'hba995023),
	.w2(32'hbba7d1b2),
	.w3(32'hbb333c59),
	.w4(32'hbb7bc9e1),
	.w5(32'hbbf6c071),
	.w6(32'h3b0e83f0),
	.w7(32'hbb30e45c),
	.w8(32'h3b1b6859),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb32c0d7),
	.w1(32'hbb258c28),
	.w2(32'hbb02bcc5),
	.w3(32'hbb0a0180),
	.w4(32'hbbe323af),
	.w5(32'hbb81f203),
	.w6(32'h3b738d4c),
	.w7(32'hbb36518b),
	.w8(32'hbaf816a9),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbf3e46),
	.w1(32'hb9b90672),
	.w2(32'hbbda499a),
	.w3(32'hbadbeb23),
	.w4(32'h3b941dbe),
	.w5(32'h39548714),
	.w6(32'hbbddafe9),
	.w7(32'h39c5e1e9),
	.w8(32'hbc20813b),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc01cb90),
	.w1(32'h3b5be012),
	.w2(32'h3c364e8a),
	.w3(32'hbc22a83a),
	.w4(32'h3b62c4de),
	.w5(32'h3c5bd734),
	.w6(32'hbc2431c5),
	.w7(32'hbaa1bcbe),
	.w8(32'h3c31f6e2),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0aae89),
	.w1(32'h3902f616),
	.w2(32'h3b22a1a7),
	.w3(32'h3c16bf00),
	.w4(32'hbc49b049),
	.w5(32'hbbeaae65),
	.w6(32'hba56bc80),
	.w7(32'hbc585910),
	.w8(32'hbc1a978d),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd15fa8),
	.w1(32'h3b5350b5),
	.w2(32'hba242dbf),
	.w3(32'hbc1fb71c),
	.w4(32'h3ba86f4b),
	.w5(32'h3bafaac7),
	.w6(32'hbb3f15a5),
	.w7(32'h3bfdc8c2),
	.w8(32'h3a80025e),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0b96f3),
	.w1(32'hbb28c3e0),
	.w2(32'hbb505c23),
	.w3(32'hb8804a53),
	.w4(32'hbb4d909d),
	.w5(32'hbbcc77e3),
	.w6(32'hba94feee),
	.w7(32'hba024f86),
	.w8(32'h3b9c8a70),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb194ea3),
	.w1(32'h3abd86cc),
	.w2(32'h3a85c43f),
	.w3(32'hbb00c595),
	.w4(32'hba90f5f4),
	.w5(32'hbc33b878),
	.w6(32'hbb17decd),
	.w7(32'hba065bc1),
	.w8(32'h3bada288),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b17a6d8),
	.w1(32'h3a153d12),
	.w2(32'hbb04240d),
	.w3(32'hbbaac220),
	.w4(32'h3ab1bbfe),
	.w5(32'hbc1ea202),
	.w6(32'hbb5c05eb),
	.w7(32'hbb3dc6c5),
	.w8(32'hbb2285b9),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3afec2),
	.w1(32'hbb933bac),
	.w2(32'hbba3bfdc),
	.w3(32'hbac91636),
	.w4(32'hbb954fb2),
	.w5(32'hbb97650b),
	.w6(32'h3b0b14a6),
	.w7(32'hbbe5fcde),
	.w8(32'hbc32c33e),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f753bf),
	.w1(32'h3b09036b),
	.w2(32'h3a833144),
	.w3(32'hbb2b6e63),
	.w4(32'h3bfd9135),
	.w5(32'hbab9e90a),
	.w6(32'hbb25a7e8),
	.w7(32'h3a979976),
	.w8(32'hbbdf8dc0),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule