module layer_8_featuremap_105(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a78f51f),
	.w1(32'hbc19996a),
	.w2(32'hbb389b84),
	.w3(32'hbb84d780),
	.w4(32'hbc261e71),
	.w5(32'hbb8e3ca5),
	.w6(32'h3ac024d0),
	.w7(32'h3b37d619),
	.w8(32'hbcff0207),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3d47e4),
	.w1(32'h3b769d7c),
	.w2(32'hbba13ab3),
	.w3(32'h3a597058),
	.w4(32'h3b550fa5),
	.w5(32'hbb3875ad),
	.w6(32'h3c1927b6),
	.w7(32'h3c81b034),
	.w8(32'hbab1fcfa),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0af97a),
	.w1(32'h3c4104ec),
	.w2(32'hbaa5a9f1),
	.w3(32'hbbeeb2f4),
	.w4(32'h38d21ac6),
	.w5(32'hbbc00924),
	.w6(32'hbb46fbfa),
	.w7(32'h3c30b073),
	.w8(32'hbc161480),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9373f6),
	.w1(32'hbcc61b2f),
	.w2(32'h3c5ce75b),
	.w3(32'h3b445f24),
	.w4(32'hbb9e55ff),
	.w5(32'h3787030c),
	.w6(32'hbc0b4e69),
	.w7(32'hbcf7f807),
	.w8(32'h3c887fef),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc12228b),
	.w1(32'hbb0d66f9),
	.w2(32'h3c0c46bb),
	.w3(32'hbc4c6567),
	.w4(32'h3c879043),
	.w5(32'hbc81daf6),
	.w6(32'hbc5653e7),
	.w7(32'hbb939109),
	.w8(32'h3a8f0036),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8cb901),
	.w1(32'h3c20d8d9),
	.w2(32'h3b8a7221),
	.w3(32'h3c192db0),
	.w4(32'h3c310a02),
	.w5(32'hbce2d171),
	.w6(32'h3bca1a17),
	.w7(32'h3c8eadd2),
	.w8(32'h3d8ff069),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb2fb84),
	.w1(32'h3c43ee99),
	.w2(32'hbc5e5a0d),
	.w3(32'hbc19f710),
	.w4(32'hbc5db17f),
	.w5(32'hbca2afc7),
	.w6(32'hbc0cad5d),
	.w7(32'hbcbe2aa4),
	.w8(32'h3c1e0132),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc59ec05),
	.w1(32'h3ba5b975),
	.w2(32'h3c460ba3),
	.w3(32'hbca5afcc),
	.w4(32'hbae36787),
	.w5(32'hbc54cf51),
	.w6(32'hbc9072ac),
	.w7(32'hbc486e7a),
	.w8(32'h3c2b7233),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9f6db3),
	.w1(32'hbb2f4d87),
	.w2(32'h3bcc99a3),
	.w3(32'hbb70b93b),
	.w4(32'hbbba2a9e),
	.w5(32'hbaf2d641),
	.w6(32'hbce753f3),
	.w7(32'hbc703f79),
	.w8(32'hba5e2cb2),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3cf0e2),
	.w1(32'h3b6be818),
	.w2(32'h3b055a12),
	.w3(32'hbb1dd855),
	.w4(32'hbbab985e),
	.w5(32'hbc8d24ee),
	.w6(32'hbbda39c1),
	.w7(32'h3c7c3092),
	.w8(32'h3a987616),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3ce5e1),
	.w1(32'hbcb2c02e),
	.w2(32'hbca8496f),
	.w3(32'hbbbe01f5),
	.w4(32'hbca91f67),
	.w5(32'hbb08d6c6),
	.w6(32'hbc557775),
	.w7(32'hbc925c33),
	.w8(32'hbc98bccc),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe31f4d),
	.w1(32'hbb31eaa6),
	.w2(32'h3c1f5a5b),
	.w3(32'hbbf7e7fe),
	.w4(32'hbbc39d36),
	.w5(32'h3c1d2b65),
	.w6(32'hbb3d82a3),
	.w7(32'hbbd27f38),
	.w8(32'h3d0e0d36),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb968fa),
	.w1(32'h3ccff6ad),
	.w2(32'h3c4c79d9),
	.w3(32'hbc826780),
	.w4(32'h3ae998ab),
	.w5(32'h3ae5584a),
	.w6(32'hbba4b275),
	.w7(32'h3c0add5f),
	.w8(32'h3c3e00f5),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4ea032),
	.w1(32'hbbb0f83b),
	.w2(32'hbab57f92),
	.w3(32'h3c24fb6f),
	.w4(32'h3b28ed1c),
	.w5(32'hbbfc652f),
	.w6(32'hbbc972c4),
	.w7(32'hbafb1aa8),
	.w8(32'hbab9558b),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd96a19),
	.w1(32'hbb48e1f8),
	.w2(32'hb98b726b),
	.w3(32'h3ae9c0c6),
	.w4(32'hbb04b586),
	.w5(32'hbc3c6d47),
	.w6(32'hbba9afc5),
	.w7(32'hbb364b9a),
	.w8(32'hbbd5e28b),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe36ee8),
	.w1(32'hbb1c4fbb),
	.w2(32'hbb44ecec),
	.w3(32'hba13b673),
	.w4(32'hbc09ed94),
	.w5(32'h3b8739f8),
	.w6(32'hbb3b77b0),
	.w7(32'hbad8a776),
	.w8(32'hbc69608f),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb836962),
	.w1(32'h3c823e5f),
	.w2(32'hbb99101d),
	.w3(32'hba510f1d),
	.w4(32'hbaa572cd),
	.w5(32'hbc4d6e38),
	.w6(32'hbc086de5),
	.w7(32'hbbd9a66b),
	.w8(32'hbc4fca09),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb917ad24),
	.w1(32'h3c4384cf),
	.w2(32'hbc176c75),
	.w3(32'hbc816f2b),
	.w4(32'hbc7b35a7),
	.w5(32'h3b82bf54),
	.w6(32'h3ad5f4f9),
	.w7(32'hbbed2476),
	.w8(32'hbcf53f40),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c299f51),
	.w1(32'hbc0f8308),
	.w2(32'hb8183816),
	.w3(32'hbd040526),
	.w4(32'hbc90ff01),
	.w5(32'h3b1d4509),
	.w6(32'h3c9baf39),
	.w7(32'hbcdb253d),
	.w8(32'hbce95389),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc87cd02),
	.w1(32'hbc6b632e),
	.w2(32'h3bbb8a99),
	.w3(32'hbc95673c),
	.w4(32'hbc40d1a5),
	.w5(32'hbd00ee46),
	.w6(32'h3b8e85a3),
	.w7(32'hbcaa9948),
	.w8(32'h3cb14e4c),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b67f7f8),
	.w1(32'hbc0bd19a),
	.w2(32'hbc117e75),
	.w3(32'h3c5f6b70),
	.w4(32'hbb9d1141),
	.w5(32'h3b9740b9),
	.w6(32'h3d0d90e9),
	.w7(32'hbbf33309),
	.w8(32'hbafc960f),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf2d8f5),
	.w1(32'h3c89734b),
	.w2(32'hbab5e4cf),
	.w3(32'h3ac69121),
	.w4(32'hbb7edf30),
	.w5(32'h3b8d55ab),
	.w6(32'hbc900065),
	.w7(32'h3b8726bc),
	.w8(32'h3d01724d),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc3e92e),
	.w1(32'hbc1816f1),
	.w2(32'hbaefe352),
	.w3(32'hbc1525ec),
	.w4(32'hbd07f867),
	.w5(32'h3c4eddcb),
	.w6(32'hbc31bd42),
	.w7(32'hbca17352),
	.w8(32'h3cad7d30),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b810992),
	.w1(32'h3b874393),
	.w2(32'hbb8f431b),
	.w3(32'h3baacc81),
	.w4(32'h3bd6d120),
	.w5(32'hbbec1dfa),
	.w6(32'hbbab8cdd),
	.w7(32'h3b85fdda),
	.w8(32'hbb479d43),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc202f23),
	.w1(32'hbb76f745),
	.w2(32'h3be3a740),
	.w3(32'h3b1ff964),
	.w4(32'hbb912857),
	.w5(32'h3bbf9b1e),
	.w6(32'hbb0cad3d),
	.w7(32'h3a2e9a83),
	.w8(32'h3c2fbb14),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c134c8f),
	.w1(32'h3a889af6),
	.w2(32'h3ba18a01),
	.w3(32'hbb9a0c15),
	.w4(32'hbc2890ca),
	.w5(32'hbc47e316),
	.w6(32'h3c316837),
	.w7(32'hb94bfd54),
	.w8(32'hbbf939ab),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8da7a5),
	.w1(32'h3d14d754),
	.w2(32'h3c36c819),
	.w3(32'h3be5221d),
	.w4(32'h3c08cd84),
	.w5(32'hbb86d41f),
	.w6(32'hbbfa173b),
	.w7(32'hbc18dfcd),
	.w8(32'hbcb514dd),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d89b09a),
	.w1(32'h3ca38439),
	.w2(32'hbcaefe3c),
	.w3(32'h3db54dc5),
	.w4(32'h3cded935),
	.w5(32'h3ca338d6),
	.w6(32'h3dc131d3),
	.w7(32'hbcdd2fae),
	.w8(32'hbd05bb47),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0e95bd),
	.w1(32'h3cb5763e),
	.w2(32'h3aef5366),
	.w3(32'h3c47395b),
	.w4(32'hbbb4d04d),
	.w5(32'h3b1163c0),
	.w6(32'h3c9a991d),
	.w7(32'h3bf1185e),
	.w8(32'h3cc6a785),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd8bf3f),
	.w1(32'hbc385a9e),
	.w2(32'h3b937efd),
	.w3(32'h3c21db6c),
	.w4(32'h3b92610a),
	.w5(32'h3c3fc951),
	.w6(32'h3b25cd60),
	.w7(32'h3b2ef24c),
	.w8(32'h3c51d985),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb06be5),
	.w1(32'h3c9115b9),
	.w2(32'h3ac0b741),
	.w3(32'h3a6f15b8),
	.w4(32'hbb531132),
	.w5(32'hbb5dba75),
	.w6(32'hbc3ca5e8),
	.w7(32'hbb93c5b8),
	.w8(32'hbaf35a7e),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabb6d84),
	.w1(32'hbb87a7b6),
	.w2(32'hbc46c882),
	.w3(32'h3bddf0a7),
	.w4(32'hbc9c0b52),
	.w5(32'hbc5e2b69),
	.w6(32'h3a7fd397),
	.w7(32'hbc8a821b),
	.w8(32'hbbd6866b),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd5dc0c),
	.w1(32'h3d061a07),
	.w2(32'h3cd05ef1),
	.w3(32'hbbd2467f),
	.w4(32'h3bd33293),
	.w5(32'h3cdbba10),
	.w6(32'hbc0ac437),
	.w7(32'h3ce137ec),
	.w8(32'h3d83743d),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf99a03),
	.w1(32'hbd1d2360),
	.w2(32'hba701e55),
	.w3(32'h3a9d3028),
	.w4(32'h3b8073a8),
	.w5(32'h3a8f71a3),
	.w6(32'hbd184741),
	.w7(32'hbbb59828),
	.w8(32'hbcab4421),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6d8f9b),
	.w1(32'h3cc5d079),
	.w2(32'h3bf929b2),
	.w3(32'hbc08cd1f),
	.w4(32'h3c0be34e),
	.w5(32'h3bf2398a),
	.w6(32'h3d140003),
	.w7(32'h3c98896e),
	.w8(32'h3c486d8a),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba1281c),
	.w1(32'hbbc0c6b9),
	.w2(32'h3bf4b392),
	.w3(32'hba6e9bf4),
	.w4(32'hba57cc96),
	.w5(32'h3cc19412),
	.w6(32'hbbf5caf7),
	.w7(32'h3cffc2d8),
	.w8(32'h3d28bfc1),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba95dc8),
	.w1(32'hbd536875),
	.w2(32'h3b40fa05),
	.w3(32'h3c329dbe),
	.w4(32'hbbccfc60),
	.w5(32'h3ba64ada),
	.w6(32'hbd535a6b),
	.w7(32'h3b91fdd6),
	.w8(32'h3c9f1775),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc0983e),
	.w1(32'hbc67adf7),
	.w2(32'hbb88fcdb),
	.w3(32'h3b001cb3),
	.w4(32'hbbbf7d11),
	.w5(32'hbbff6827),
	.w6(32'h3b30bd1f),
	.w7(32'hbb869f95),
	.w8(32'hbc1ffa14),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab80603),
	.w1(32'h3ca35d79),
	.w2(32'hbb5d2d9f),
	.w3(32'h3c11f391),
	.w4(32'hbbffdc6f),
	.w5(32'hbc597135),
	.w6(32'h3c4751a1),
	.w7(32'hbcbd1f47),
	.w8(32'hbc7b5d34),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8548ba),
	.w1(32'h3ccaf3fa),
	.w2(32'h3c6bd8c5),
	.w3(32'hbbf5b42e),
	.w4(32'hbb6d2a95),
	.w5(32'h3b712e84),
	.w6(32'h3ced1f9c),
	.w7(32'h3a3be669),
	.w8(32'h3b867332),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b12a93c),
	.w1(32'hbc3cc262),
	.w2(32'h3c147df9),
	.w3(32'hbd25fdb9),
	.w4(32'hbcd7d723),
	.w5(32'hbbb185ed),
	.w6(32'hbc9f6129),
	.w7(32'hbc46a301),
	.w8(32'hbb9e1607),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca04c53),
	.w1(32'h3ccbed25),
	.w2(32'h3c1f38fb),
	.w3(32'hba8d106b),
	.w4(32'hbbad048d),
	.w5(32'h3c5be4cb),
	.w6(32'h3c949e8d),
	.w7(32'h3ae35f66),
	.w8(32'hbb32b609),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb1d4f9),
	.w1(32'hba994d25),
	.w2(32'h3b41dc30),
	.w3(32'hbc744a3a),
	.w4(32'h3be616d1),
	.w5(32'h3b878e6a),
	.w6(32'h3cac6c9e),
	.w7(32'h3c8a066f),
	.w8(32'h3d3a66c2),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1d64b3),
	.w1(32'hbcd8b88c),
	.w2(32'h3c238f32),
	.w3(32'h3c462162),
	.w4(32'hbbb1340d),
	.w5(32'hba592f20),
	.w6(32'hbbd8910e),
	.w7(32'hbb3c2f2a),
	.w8(32'h3c038fc6),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba85755b),
	.w1(32'hbc88711e),
	.w2(32'hbc3a1d13),
	.w3(32'h3b29f7e3),
	.w4(32'hbc6f73ee),
	.w5(32'hbb5a3c70),
	.w6(32'hbc6744ec),
	.w7(32'hbc1f7557),
	.w8(32'hbca1999e),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8ba597),
	.w1(32'h3cae7320),
	.w2(32'h3bfd5f9b),
	.w3(32'h3c4d509c),
	.w4(32'h3b933a2a),
	.w5(32'h3babc22e),
	.w6(32'h3bac2578),
	.w7(32'h3bb18714),
	.w8(32'h3d3559f8),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b21640c),
	.w1(32'hbc89d13e),
	.w2(32'h3c99b52f),
	.w3(32'hbb6c34cf),
	.w4(32'hbb289c17),
	.w5(32'hb9e4eaaf),
	.w6(32'hbcf5ef4f),
	.w7(32'h3cd53600),
	.w8(32'h3c17dced),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b71fa12),
	.w1(32'hbc882f74),
	.w2(32'h3985151c),
	.w3(32'h3bb13d93),
	.w4(32'hbaa3829d),
	.w5(32'h3c2e9c0b),
	.w6(32'hba773cb0),
	.w7(32'hbbe16fb0),
	.w8(32'h3cb3ec87),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1eae18),
	.w1(32'hbc9c012f),
	.w2(32'hbc96005c),
	.w3(32'h3b4edefd),
	.w4(32'hbbb5ee57),
	.w5(32'hbb75e4ff),
	.w6(32'hbcd84462),
	.w7(32'hbb9ee531),
	.w8(32'hbd451a38),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3caf7f3c),
	.w1(32'h3c506abc),
	.w2(32'hbd17bc61),
	.w3(32'hbcd40ed4),
	.w4(32'hbd49efb9),
	.w5(32'hbd32ac9c),
	.w6(32'h3cd06dd4),
	.w7(32'hbd6959f7),
	.w8(32'hbcfc1593),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cdd1ca5),
	.w1(32'h3d64f87b),
	.w2(32'hbb8af641),
	.w3(32'hbc4bbc50),
	.w4(32'h3b51b7d8),
	.w5(32'hbbeeaca6),
	.w6(32'h3d575251),
	.w7(32'h3c3ccf0d),
	.w8(32'hbb8bfdf2),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd0ab3d),
	.w1(32'h3c289d53),
	.w2(32'h3c60fb2c),
	.w3(32'hbc05144a),
	.w4(32'hbca9b5d0),
	.w5(32'h3a9b2d0b),
	.w6(32'hbc8fb44d),
	.w7(32'hbce3903e),
	.w8(32'h3ccd42df),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf180b9),
	.w1(32'h3c9e7dc3),
	.w2(32'hbc967277),
	.w3(32'hbbfb8b63),
	.w4(32'hba8f9d34),
	.w5(32'hbc580903),
	.w6(32'hba3ebed4),
	.w7(32'hbc5f0844),
	.w8(32'hbcce02c8),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb61aa3),
	.w1(32'hbc07be3f),
	.w2(32'h3b2c35d9),
	.w3(32'hbd15ab12),
	.w4(32'hbc688bf8),
	.w5(32'hbc46fe49),
	.w6(32'hbc7176cf),
	.w7(32'hbc0ac2d1),
	.w8(32'h3a7662b9),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaff9bc4),
	.w1(32'hbc04fad1),
	.w2(32'h3c52ffa3),
	.w3(32'h3c006656),
	.w4(32'hbc2ae000),
	.w5(32'h3bc0adbc),
	.w6(32'hbbb3d427),
	.w7(32'h3c74378a),
	.w8(32'h3be74101),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc53561d),
	.w1(32'hbb91af28),
	.w2(32'hbbc90db9),
	.w3(32'hbb5c066e),
	.w4(32'hbcec6d46),
	.w5(32'hbcf8a7e0),
	.w6(32'hbc8081cb),
	.w7(32'hbd04d94c),
	.w8(32'hbc30092f),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7f2ffb),
	.w1(32'h3c004838),
	.w2(32'hbc1bbebf),
	.w3(32'h3c805057),
	.w4(32'h3bba6f73),
	.w5(32'hb9d69ba0),
	.w6(32'h3c88e1ce),
	.w7(32'hbaf1984e),
	.w8(32'hbc69f6a3),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc496f74),
	.w1(32'h3acb35d7),
	.w2(32'h3c488a35),
	.w3(32'hbc80c9ba),
	.w4(32'h3a89359b),
	.w5(32'h3c81b105),
	.w6(32'hbcb7880d),
	.w7(32'hbbd0e2b7),
	.w8(32'h3c6f234d),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc192e15),
	.w1(32'h3b3a223b),
	.w2(32'h3c06987a),
	.w3(32'h3c87d695),
	.w4(32'h39a7cd12),
	.w5(32'h3b5858b3),
	.w6(32'h3c2258e2),
	.w7(32'hba353ef7),
	.w8(32'h3c216cf5),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbea9c98),
	.w1(32'hbc572e00),
	.w2(32'hbbc13ec2),
	.w3(32'h3b9d01f5),
	.w4(32'hbbe1dfd4),
	.w5(32'hbc2b63eb),
	.w6(32'hbbfaae32),
	.w7(32'hbc4661cd),
	.w8(32'hbc95865b),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8e7078),
	.w1(32'h3c6d87dc),
	.w2(32'hbc70e89f),
	.w3(32'h3bb8e6e5),
	.w4(32'hbbe783aa),
	.w5(32'hbc8c7c5b),
	.w6(32'h3c2faffe),
	.w7(32'hbc97adca),
	.w8(32'h3c55a2d6),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8bbac6),
	.w1(32'h3c071a8e),
	.w2(32'hbb681023),
	.w3(32'h3cafaf75),
	.w4(32'h3ac3b21f),
	.w5(32'hbb9652d3),
	.w6(32'h3c803be7),
	.w7(32'h3b0c61e1),
	.w8(32'hba179cdf),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca0b796),
	.w1(32'hbc7cb942),
	.w2(32'h3a7e6447),
	.w3(32'hbc375569),
	.w4(32'hbcd2fd1f),
	.w5(32'hbcf02ee9),
	.w6(32'hbb7bc0bf),
	.w7(32'hbc8c295c),
	.w8(32'hbce74095),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb9f5e3),
	.w1(32'hbc3a216c),
	.w2(32'h3bb6c258),
	.w3(32'hbc324a3d),
	.w4(32'h3adeb3b4),
	.w5(32'h3b153d40),
	.w6(32'hbca055b0),
	.w7(32'hbc29db2c),
	.w8(32'hbc1ded5e),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa83a78),
	.w1(32'h3c741d2b),
	.w2(32'h3af18f20),
	.w3(32'h3bb23a1a),
	.w4(32'hb8d76c22),
	.w5(32'h3c6f4135),
	.w6(32'h3b5e42f3),
	.w7(32'h3c55d164),
	.w8(32'h3c3dc4d3),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc075162),
	.w1(32'hbc22d637),
	.w2(32'h39667f37),
	.w3(32'hbb524e3c),
	.w4(32'h3bde12fc),
	.w5(32'h3acdf318),
	.w6(32'hbc8ac587),
	.w7(32'h3be5efc8),
	.w8(32'h3bc4b426),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbba7be8),
	.w1(32'h3aef0c46),
	.w2(32'h3b904297),
	.w3(32'hbc0399bf),
	.w4(32'h3b8b661e),
	.w5(32'h3c063171),
	.w6(32'h3b2af133),
	.w7(32'h3c162dfc),
	.w8(32'hbb7da7b4),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc17e84a),
	.w1(32'h3cbd63c9),
	.w2(32'h3ca354a7),
	.w3(32'hbb193b8b),
	.w4(32'h3aee7a7f),
	.w5(32'h3c03f357),
	.w6(32'h3cdda6fa),
	.w7(32'hba3fc04a),
	.w8(32'hbadd5448),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca0a8e1),
	.w1(32'h3c062403),
	.w2(32'h3bab5eca),
	.w3(32'hbcd42569),
	.w4(32'hbab437a4),
	.w5(32'hbc1bc945),
	.w6(32'hbcecf2ff),
	.w7(32'hbc32baf3),
	.w8(32'hbcd43e33),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6d5eb3),
	.w1(32'hbba10300),
	.w2(32'hbd0742f0),
	.w3(32'h3c2ad0ab),
	.w4(32'hbc56cda7),
	.w5(32'hbc8e1965),
	.w6(32'h3d4a0bf8),
	.w7(32'hbccf1186),
	.w8(32'hbcd39fdb),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc2bb41),
	.w1(32'hbbc89b3b),
	.w2(32'hbc2154be),
	.w3(32'hbc8144f3),
	.w4(32'hbc3ae5ed),
	.w5(32'h3bbe618c),
	.w6(32'h3a5471c3),
	.w7(32'hbb97d0b6),
	.w8(32'hbc1d420d),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb88e764),
	.w1(32'hbb9edd75),
	.w2(32'hbba0e82d),
	.w3(32'hbce5493e),
	.w4(32'hbaf66521),
	.w5(32'hbc98b604),
	.w6(32'h3b0cecd2),
	.w7(32'h399a008c),
	.w8(32'hbcf894d9),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d1fbd02),
	.w1(32'hbc03633c),
	.w2(32'h3beace26),
	.w3(32'h3cdd7a15),
	.w4(32'hbbad61eb),
	.w5(32'hbb959ea3),
	.w6(32'h3d2cff92),
	.w7(32'hbc45fbd9),
	.w8(32'h3bee0a01),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c816b4a),
	.w1(32'h3c75b9c5),
	.w2(32'h3b97e191),
	.w3(32'hbc98b32e),
	.w4(32'hbb95b8d5),
	.w5(32'hbb43b69c),
	.w6(32'hbc0fc4af),
	.w7(32'hbbf78d34),
	.w8(32'hbb7c9203),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb558b48),
	.w1(32'hbb59c069),
	.w2(32'h3c290897),
	.w3(32'hbc4e1753),
	.w4(32'hbc781a2f),
	.w5(32'hbbfc393b),
	.w6(32'hbba28b09),
	.w7(32'hbc07a990),
	.w8(32'hbc9a5b46),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b25386),
	.w1(32'h3c9b2502),
	.w2(32'h3bad26f3),
	.w3(32'hbb4e697b),
	.w4(32'h3c4d60e0),
	.w5(32'hbc52eab4),
	.w6(32'h3bb08103),
	.w7(32'hbaf0690e),
	.w8(32'h3c7e2ac2),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d3ebfb5),
	.w1(32'hbc327cbd),
	.w2(32'h3b99e468),
	.w3(32'h3cb24d1b),
	.w4(32'h3a42aab7),
	.w5(32'h3b4a4fc0),
	.w6(32'h3c1db152),
	.w7(32'hbae7d36c),
	.w8(32'h3bef1bae),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe26b47),
	.w1(32'hbbb7fa94),
	.w2(32'h3b756141),
	.w3(32'hbb72d8f6),
	.w4(32'hb9d1136a),
	.w5(32'h3aab2724),
	.w6(32'hba0e8e47),
	.w7(32'hbc1cf158),
	.w8(32'hbb94ebdf),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b166812),
	.w1(32'h3c022b16),
	.w2(32'h3c1fd9fb),
	.w3(32'hbc1c7559),
	.w4(32'hbb835b02),
	.w5(32'hbb068bf9),
	.w6(32'h3a8e9aaf),
	.w7(32'hbc24b0cf),
	.w8(32'hbba911bb),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba84123d),
	.w1(32'h3bfe9fb2),
	.w2(32'hbbe0e988),
	.w3(32'h3b0dc0ea),
	.w4(32'h3b90f520),
	.w5(32'hb927e205),
	.w6(32'h3b92b47f),
	.w7(32'hbafa1ff6),
	.w8(32'hbc8c3c20),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdb0feb),
	.w1(32'hbbf1de74),
	.w2(32'hbbac6695),
	.w3(32'hbc221dc6),
	.w4(32'hbc438760),
	.w5(32'hbb926b01),
	.w6(32'h3c1579a7),
	.w7(32'hbbd78545),
	.w8(32'hbc6b7192),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc373a40),
	.w1(32'hbc45fd6c),
	.w2(32'hbb32d663),
	.w3(32'hb9988330),
	.w4(32'h3cc49e47),
	.w5(32'hbc373b9c),
	.w6(32'h3a57e4c0),
	.w7(32'hbc61b420),
	.w8(32'h3c77eda8),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc361e1a),
	.w1(32'hbcc9efcf),
	.w2(32'hbaad2977),
	.w3(32'hbb1c7a8e),
	.w4(32'hbca4d7e6),
	.w5(32'hbba01c30),
	.w6(32'hbc835829),
	.w7(32'hbc39a266),
	.w8(32'hbca67705),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc85cad0),
	.w1(32'hbcbb29a3),
	.w2(32'h3b93da0e),
	.w3(32'hbcf87406),
	.w4(32'hbc633cd3),
	.w5(32'hbc2d8cbe),
	.w6(32'hbd0fd84d),
	.w7(32'h3bb4d19d),
	.w8(32'hbb7b79bf),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4752ce),
	.w1(32'hbcb1610f),
	.w2(32'hbc8fb3a4),
	.w3(32'hbc4b5a6c),
	.w4(32'hbd2c91b1),
	.w5(32'h3cf9081d),
	.w6(32'hba76430a),
	.w7(32'hbbde28c4),
	.w8(32'hbd721687),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb372564),
	.w1(32'hbc50be01),
	.w2(32'hbc12d623),
	.w3(32'hbd0e88fe),
	.w4(32'hbc198c20),
	.w5(32'hbc06d68a),
	.w6(32'h3d1369fe),
	.w7(32'h3a2d7eb9),
	.w8(32'hbcb06524),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c298b3f),
	.w1(32'h3a8a4f65),
	.w2(32'hbb92b93a),
	.w3(32'hbb29db7b),
	.w4(32'h3b875607),
	.w5(32'hbaa04314),
	.w6(32'hbc1315a4),
	.w7(32'h3ae1b995),
	.w8(32'hbd1034fd),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8780cd),
	.w1(32'hb9c7819a),
	.w2(32'h3c0828b9),
	.w3(32'h3ad6bb73),
	.w4(32'h3c7dbf63),
	.w5(32'hbb66c77c),
	.w6(32'h3c7524be),
	.w7(32'h3acd6bbb),
	.w8(32'h3c0d4b75),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b68c0df),
	.w1(32'h393c8e9f),
	.w2(32'hba9e482b),
	.w3(32'hbb4b431a),
	.w4(32'h3b0fb2ab),
	.w5(32'hbb1f065b),
	.w6(32'hbb5d4959),
	.w7(32'h3b876fe3),
	.w8(32'hbbfcafa1),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5a7220),
	.w1(32'hbbb22618),
	.w2(32'hbc32cb75),
	.w3(32'hbc30d931),
	.w4(32'hbcae2eda),
	.w5(32'h3d09a801),
	.w6(32'h3bfe96e3),
	.w7(32'h3c664949),
	.w8(32'hbdbdecdd),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac14ab3),
	.w1(32'h3c15924b),
	.w2(32'hbb0a4a1d),
	.w3(32'hbcd49909),
	.w4(32'h3c0c5f24),
	.w5(32'hbc7e6a96),
	.w6(32'h3d37bd82),
	.w7(32'hbbd4ce02),
	.w8(32'hbc11fa6b),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c20f05f),
	.w1(32'hbc63d92e),
	.w2(32'h3c37fc93),
	.w3(32'h3b130d4e),
	.w4(32'hbbb9125e),
	.w5(32'hba1d4a02),
	.w6(32'hba8b16a6),
	.w7(32'hba1db808),
	.w8(32'hbbd42630),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc882c54),
	.w1(32'h3b8e9d70),
	.w2(32'hbc1ad458),
	.w3(32'hbbacb0ac),
	.w4(32'h3a4663c9),
	.w5(32'hbbb50124),
	.w6(32'hbbc2aec8),
	.w7(32'h3b599583),
	.w8(32'hbba1c102),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2a6d9c),
	.w1(32'hba0b8716),
	.w2(32'h3c350388),
	.w3(32'hbbb5efa7),
	.w4(32'h3b6cd5f5),
	.w5(32'h3c2c8913),
	.w6(32'h3b9f2504),
	.w7(32'hbcc7952c),
	.w8(32'h3d6d3aad),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd2e772f),
	.w1(32'h3c7144b2),
	.w2(32'h3baae102),
	.w3(32'hbc4dbe48),
	.w4(32'h3b108512),
	.w5(32'hba369a1b),
	.w6(32'hbca2e904),
	.w7(32'h392ecdc3),
	.w8(32'hbb98b39a),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba4622d),
	.w1(32'hb9e60686),
	.w2(32'h3b89ccf4),
	.w3(32'h3bf59221),
	.w4(32'hbbba9034),
	.w5(32'hbbd77294),
	.w6(32'h3a668563),
	.w7(32'hbc5f59d5),
	.w8(32'h3c346a64),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc69aa0),
	.w1(32'h3ba92bd5),
	.w2(32'h3ad9751e),
	.w3(32'hbc81f57c),
	.w4(32'hbca4dd41),
	.w5(32'h3cbe4e9d),
	.w6(32'hbcb11ab6),
	.w7(32'hbcb0f6dc),
	.w8(32'h3a705fbf),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3faa10),
	.w1(32'hbb1fb81c),
	.w2(32'hba5b56f1),
	.w3(32'hbc06c3b7),
	.w4(32'h3c48219b),
	.w5(32'h3b807924),
	.w6(32'hbc1ab765),
	.w7(32'hbc8cf7b3),
	.w8(32'h3c162959),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca24f58),
	.w1(32'hba3a348c),
	.w2(32'h3a70aa02),
	.w3(32'hbc911095),
	.w4(32'hbb126c9d),
	.w5(32'h3bb3daab),
	.w6(32'h3c345248),
	.w7(32'h3b3481d9),
	.w8(32'hbbc86ac1),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a83605d),
	.w1(32'h3b4e63f8),
	.w2(32'h3c4b547f),
	.w3(32'h3bb466b7),
	.w4(32'hbc00024d),
	.w5(32'h3c123e90),
	.w6(32'h3b988a5b),
	.w7(32'hbbc52c2c),
	.w8(32'h3c94b79e),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc29b0f1),
	.w1(32'hbc0f2abe),
	.w2(32'h3c4e57fc),
	.w3(32'h3ba9d488),
	.w4(32'h3b987524),
	.w5(32'h3be145f3),
	.w6(32'hbbf1c93c),
	.w7(32'h3c522256),
	.w8(32'hbc890489),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc73196c),
	.w1(32'h3be23029),
	.w2(32'hbc08c662),
	.w3(32'hbb1bcc33),
	.w4(32'h3c2102c4),
	.w5(32'hbc32a564),
	.w6(32'hbaaa6473),
	.w7(32'h3b3bf725),
	.w8(32'h3c5c1725),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6d61fd),
	.w1(32'h3c4d99f2),
	.w2(32'h3b1844b4),
	.w3(32'hb9d3bbb0),
	.w4(32'hbb81ca1f),
	.w5(32'h3bf60a03),
	.w6(32'h3bf8feab),
	.w7(32'hbbc2ed0c),
	.w8(32'hbc643627),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6a08d1),
	.w1(32'hbba92399),
	.w2(32'hbbe28c82),
	.w3(32'h3b92d320),
	.w4(32'h3bb732f4),
	.w5(32'hb999a048),
	.w6(32'hbba51629),
	.w7(32'h3ba71c5f),
	.w8(32'hba8d4e95),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba024dfe),
	.w1(32'h3b098d8a),
	.w2(32'hbc29b459),
	.w3(32'h3c1f965a),
	.w4(32'hbb83ba88),
	.w5(32'hbc3cb2dd),
	.w6(32'hbb37aa82),
	.w7(32'hbc0e1ee4),
	.w8(32'h3cc7f965),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c262feb),
	.w1(32'h39559026),
	.w2(32'hba3ea544),
	.w3(32'hbc073a67),
	.w4(32'h3ba59088),
	.w5(32'h3ba9d8a8),
	.w6(32'h3bc6b3f3),
	.w7(32'hb9337f05),
	.w8(32'hbc9ca7b0),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c53a105),
	.w1(32'hbc237a74),
	.w2(32'hbc021df0),
	.w3(32'h3c589103),
	.w4(32'h3aee70cf),
	.w5(32'hbce1d774),
	.w6(32'h3c6730b3),
	.w7(32'hbc5add9f),
	.w8(32'h3cc40681),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c53b828),
	.w1(32'h3ad6b276),
	.w2(32'h3c231471),
	.w3(32'h3c7f58c0),
	.w4(32'h3bb6f56e),
	.w5(32'h3c15d194),
	.w6(32'hbcaa9914),
	.w7(32'h3b414b66),
	.w8(32'h3c7aab78),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2b68f1),
	.w1(32'h3b5bb342),
	.w2(32'hb9d87906),
	.w3(32'h39eb6334),
	.w4(32'hbb078161),
	.w5(32'hbba35178),
	.w6(32'hba80a58e),
	.w7(32'h3c0d63e2),
	.w8(32'hbb242219),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9d76ec),
	.w1(32'hbc125fe4),
	.w2(32'h3ac031f9),
	.w3(32'hb987c636),
	.w4(32'h3c585a4b),
	.w5(32'hbd80047b),
	.w6(32'h3ba8673a),
	.w7(32'hbd0a08cc),
	.w8(32'h3d5b946a),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b40dc75),
	.w1(32'hba2d62a6),
	.w2(32'hbbb2bc91),
	.w3(32'h3d0462f3),
	.w4(32'h3a46903d),
	.w5(32'h3c4d46e0),
	.w6(32'hbd21198c),
	.w7(32'h3c3c0a8e),
	.w8(32'hbc7e648d),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f2e544),
	.w1(32'h3b99647e),
	.w2(32'h3bad9d27),
	.w3(32'hbc656ec4),
	.w4(32'h39b4ad28),
	.w5(32'h3c1984bd),
	.w6(32'h3c41d308),
	.w7(32'hbba2e9c7),
	.w8(32'hbb6737ea),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc20f04e),
	.w1(32'h3af30f28),
	.w2(32'hba47182f),
	.w3(32'hbc9831e3),
	.w4(32'h3c0630c7),
	.w5(32'hbc8cb8ed),
	.w6(32'hbc285841),
	.w7(32'hbc7c7f64),
	.w8(32'h3c152b3d),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3759ead8),
	.w1(32'hbd10cf1d),
	.w2(32'hbc404f5e),
	.w3(32'hbb0fc9cb),
	.w4(32'hbc7b954d),
	.w5(32'hbc6ae94e),
	.w6(32'h3a9e00df),
	.w7(32'hbc5b36a8),
	.w8(32'h3a9373f5),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc938fae),
	.w1(32'hbcd628c4),
	.w2(32'hbc1fbcfe),
	.w3(32'hbc52e78c),
	.w4(32'h3b2b7078),
	.w5(32'hbca8dc46),
	.w6(32'hbc7e1507),
	.w7(32'h3bed6513),
	.w8(32'h3c612531),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc812d28),
	.w1(32'hbc009dbc),
	.w2(32'hbc8a5838),
	.w3(32'hbc681daa),
	.w4(32'hbb327bfb),
	.w5(32'h3c5a957f),
	.w6(32'hba0aeff2),
	.w7(32'h3c5f97b8),
	.w8(32'hbca8ea5a),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad95f86),
	.w1(32'h3c7b0e40),
	.w2(32'h399d509b),
	.w3(32'hbc110c65),
	.w4(32'hbc6ff72d),
	.w5(32'hbc042f70),
	.w6(32'h3bd2bb17),
	.w7(32'h3af66dc4),
	.w8(32'h3d54e579),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc80e0e0),
	.w1(32'h3c68db45),
	.w2(32'h3c0e4bb0),
	.w3(32'hbc0c1bfa),
	.w4(32'hbb938f45),
	.w5(32'h3bc63f49),
	.w6(32'hbcc30782),
	.w7(32'hbbb9f8aa),
	.w8(32'h3bd6d0cf),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39632acd),
	.w1(32'h3b5d5ada),
	.w2(32'hbbca8dc8),
	.w3(32'hba29baa3),
	.w4(32'hbc0315b2),
	.w5(32'hbbe87f86),
	.w6(32'hbb0cdaf7),
	.w7(32'h3b938374),
	.w8(32'h3b7bdd8a),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a87e5),
	.w1(32'h3c11117e),
	.w2(32'h3b1a9858),
	.w3(32'h3a950ab3),
	.w4(32'hbc8b256a),
	.w5(32'hbc2c833f),
	.w6(32'hbbc856c8),
	.w7(32'hb97e5e88),
	.w8(32'h3c518489),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc099656),
	.w1(32'hbc8bae57),
	.w2(32'hbbd2335d),
	.w3(32'hbb87f3dc),
	.w4(32'h3aba876a),
	.w5(32'hbb1b2fb3),
	.w6(32'hbc7ddbb2),
	.w7(32'hbb913a16),
	.w8(32'h3b1974da),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aebd008),
	.w1(32'h3c6ea1cf),
	.w2(32'h3c16a447),
	.w3(32'hb8c6c62c),
	.w4(32'h3bc833e7),
	.w5(32'h3a1a61f0),
	.w6(32'h3b8bda8e),
	.w7(32'h3c8a1674),
	.w8(32'hbc0ef53d),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c36c05),
	.w1(32'h3b33023f),
	.w2(32'h3c15d4c0),
	.w3(32'hbb0c8e5a),
	.w4(32'h3ad3b25a),
	.w5(32'h3bd822cd),
	.w6(32'hbb4edd48),
	.w7(32'hbae7b3e0),
	.w8(32'h3c2843ae),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a867a91),
	.w1(32'h3bbdb305),
	.w2(32'hbc63891f),
	.w3(32'h3a1405fb),
	.w4(32'hbbd8077a),
	.w5(32'h3c845f28),
	.w6(32'hbb187d0f),
	.w7(32'h3d21bcac),
	.w8(32'hbdaac736),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce2b7b6),
	.w1(32'hbc43d93b),
	.w2(32'h3c312023),
	.w3(32'h3af9f100),
	.w4(32'h3b8a7c45),
	.w5(32'hbc949ddc),
	.w6(32'h3d0fb036),
	.w7(32'hbc5f98fd),
	.w8(32'h3d4ca434),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1e25d1),
	.w1(32'h3b380094),
	.w2(32'h3b94044f),
	.w3(32'h3c9c8add),
	.w4(32'h3ba5873c),
	.w5(32'h3ad3bbaf),
	.w6(32'hbbc4d017),
	.w7(32'h3b8999df),
	.w8(32'hbb56a656),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a16e781),
	.w1(32'h3bd0c7f1),
	.w2(32'hbaf3f804),
	.w3(32'hba848b99),
	.w4(32'hbacb3372),
	.w5(32'hbbd09bdf),
	.w6(32'h3b590977),
	.w7(32'h3c0b37ed),
	.w8(32'hbc5086b7),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c158369),
	.w1(32'h3b44370a),
	.w2(32'h3c34fae5),
	.w3(32'hbc327fa3),
	.w4(32'h3bcae8cc),
	.w5(32'h393fe61c),
	.w6(32'hb93c9013),
	.w7(32'hbb9ed205),
	.w8(32'h39f7987b),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule