module layer_10_featuremap_471(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb15651a),
	.w1(32'h3bd842df),
	.w2(32'hbb2323ff),
	.w3(32'hbb8d0aad),
	.w4(32'h3c4a9806),
	.w5(32'hbbeb33be),
	.w6(32'hbb8b4165),
	.w7(32'h3be39f38),
	.w8(32'h3abd1579),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb16e49d),
	.w1(32'hbaf43b5e),
	.w2(32'hba8d51ed),
	.w3(32'hbb6f35d6),
	.w4(32'hbb104f7b),
	.w5(32'h3c350702),
	.w6(32'h3adbe325),
	.w7(32'h3a428598),
	.w8(32'h3b943ff6),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb936ce14),
	.w1(32'h3a864807),
	.w2(32'hbac24c76),
	.w3(32'hbb44777a),
	.w4(32'h3c24ec1d),
	.w5(32'h3873b481),
	.w6(32'hbba97150),
	.w7(32'hbb63ce83),
	.w8(32'hbb1cafa9),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba97d106),
	.w1(32'hbb63f276),
	.w2(32'hbb4cd3eb),
	.w3(32'h3b37bcc2),
	.w4(32'hbb8dd1ea),
	.w5(32'h38af1dc3),
	.w6(32'hbb167489),
	.w7(32'hbbc02969),
	.w8(32'hbbc3167f),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf0a0a0),
	.w1(32'h3aadfd29),
	.w2(32'h3aff3d67),
	.w3(32'hbc24a7fa),
	.w4(32'h3c03f607),
	.w5(32'h3b8183b2),
	.w6(32'hbbf26d01),
	.w7(32'h3ac43e33),
	.w8(32'h3bd8e9e8),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aef651d),
	.w1(32'hbbd2678b),
	.w2(32'h3be1e76b),
	.w3(32'hb8b80814),
	.w4(32'hbc721559),
	.w5(32'h3c8df974),
	.w6(32'h3b4cd151),
	.w7(32'hbbce63cb),
	.w8(32'h3c101a0e),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc70893),
	.w1(32'hba53fded),
	.w2(32'h3bd1e101),
	.w3(32'h3ba42629),
	.w4(32'h3a3700c2),
	.w5(32'h3bea21dc),
	.w6(32'h3b692150),
	.w7(32'hb9af9d54),
	.w8(32'h3a861e41),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c233999),
	.w1(32'h3bbdd36c),
	.w2(32'h3c22bea2),
	.w3(32'h3c2f863c),
	.w4(32'h3baef2e6),
	.w5(32'h3bf24b2c),
	.w6(32'h3a38f20a),
	.w7(32'h3ae95c45),
	.w8(32'h3c149429),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b896eef),
	.w1(32'hbb97539d),
	.w2(32'hbc213e50),
	.w3(32'h3bcb6bdd),
	.w4(32'hbaf4db33),
	.w5(32'hbb55fa68),
	.w6(32'h3b6052b5),
	.w7(32'hbbb42464),
	.w8(32'hbc1278ce),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c559564),
	.w1(32'hba739bbd),
	.w2(32'h3af52350),
	.w3(32'h3c08fb80),
	.w4(32'h3b4e8673),
	.w5(32'h3b99ee24),
	.w6(32'h3ac2ba1f),
	.w7(32'h3aaf740f),
	.w8(32'h3bee05b3),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb96fe0c),
	.w1(32'hbb854991),
	.w2(32'hba53150b),
	.w3(32'hbad5451c),
	.w4(32'hbab8fac9),
	.w5(32'h3b40067c),
	.w6(32'h3bb66fce),
	.w7(32'hbb5cbb10),
	.w8(32'hba024da4),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb86ee9b),
	.w1(32'hbb648ecb),
	.w2(32'hbbce1b94),
	.w3(32'hbb831246),
	.w4(32'hba8d2fa2),
	.w5(32'hbb99ba4d),
	.w6(32'hbc329a89),
	.w7(32'hbb0a9c6b),
	.w8(32'hbc0df295),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6d6845),
	.w1(32'h3adf2eb0),
	.w2(32'hbb0a09c7),
	.w3(32'h3c16603c),
	.w4(32'h3ae57ac4),
	.w5(32'h3c930ce6),
	.w6(32'h3bbec4d9),
	.w7(32'hbb513d42),
	.w8(32'h3ac07b8a),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a071768),
	.w1(32'h3a294df2),
	.w2(32'hbb9f4187),
	.w3(32'h3abafee9),
	.w4(32'h3b3b3d4e),
	.w5(32'hbac6f945),
	.w6(32'hb921936f),
	.w7(32'hba5afd25),
	.w8(32'h380df47f),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab3cfd9),
	.w1(32'hbb5dd63b),
	.w2(32'hbb279b95),
	.w3(32'h3b8871d6),
	.w4(32'hbbc741ac),
	.w5(32'h3b146982),
	.w6(32'hba448350),
	.w7(32'hbb74b5c9),
	.w8(32'hbb75c608),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c18bab9),
	.w1(32'h3befa02e),
	.w2(32'hba6f8df9),
	.w3(32'h3bd25416),
	.w4(32'h3bf04249),
	.w5(32'h3985717d),
	.w6(32'h3be3ef96),
	.w7(32'h3be37035),
	.w8(32'h3959331a),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfc109d),
	.w1(32'h3bd59b77),
	.w2(32'h3bea0ee6),
	.w3(32'hbc1829b1),
	.w4(32'h3af9fbd5),
	.w5(32'hba80393f),
	.w6(32'hbc42c196),
	.w7(32'h3aeb895f),
	.w8(32'hbaea20cc),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8fee2d),
	.w1(32'h3be2a58d),
	.w2(32'h3c6e8642),
	.w3(32'h3c101ff3),
	.w4(32'h3b0f5047),
	.w5(32'h3a17a50c),
	.w6(32'h3bd33e3d),
	.w7(32'h3af5f2bc),
	.w8(32'hbb03b7f5),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd036dd),
	.w1(32'hba8d1cd7),
	.w2(32'h3b23c848),
	.w3(32'h3b4257aa),
	.w4(32'h3ac8094a),
	.w5(32'h3c2963f1),
	.w6(32'h3b051c01),
	.w7(32'hba9b531b),
	.w8(32'h3bab3372),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba85a71f),
	.w1(32'h3a90526f),
	.w2(32'h3ba25239),
	.w3(32'hbb984099),
	.w4(32'hbacca3fe),
	.w5(32'h3af6b076),
	.w6(32'hbb997d88),
	.w7(32'h3bb4376d),
	.w8(32'hb9b278c2),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fc432a),
	.w1(32'hbab18147),
	.w2(32'h3c0db234),
	.w3(32'hba42c30c),
	.w4(32'hbb57b834),
	.w5(32'h3c8b5e68),
	.w6(32'h3b8da875),
	.w7(32'h3a986408),
	.w8(32'h3c02c131),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b07cbd7),
	.w1(32'h39c56801),
	.w2(32'h3b8da1c2),
	.w3(32'h3ae27d27),
	.w4(32'hbc25a746),
	.w5(32'h3c3cbd16),
	.w6(32'hbab8d64e),
	.w7(32'h3a80a549),
	.w8(32'h3acded44),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b21f400),
	.w1(32'h3c2580f3),
	.w2(32'h3cb79ed4),
	.w3(32'h39d9c0a3),
	.w4(32'hbb8c2a33),
	.w5(32'h3c843148),
	.w6(32'h3b931c08),
	.w7(32'h3b99cabc),
	.w8(32'h3bbb077b),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfab189),
	.w1(32'h3c24ce85),
	.w2(32'h3bb01224),
	.w3(32'h3c81ae9a),
	.w4(32'h3baea75b),
	.w5(32'hbb331255),
	.w6(32'h3c36faf9),
	.w7(32'h3c42c85b),
	.w8(32'h3b8dfaee),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c39de27),
	.w1(32'hba0305ca),
	.w2(32'h3bc79226),
	.w3(32'h3bf3eaf9),
	.w4(32'hba596cab),
	.w5(32'h3a84a707),
	.w6(32'h3c2485b4),
	.w7(32'h37683677),
	.w8(32'hba16327a),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab1a190),
	.w1(32'hbbc046e9),
	.w2(32'h3c04aa66),
	.w3(32'h3a880ce4),
	.w4(32'hbc1f49ad),
	.w5(32'h3c526885),
	.w6(32'hb9d79a79),
	.w7(32'hbc1662ed),
	.w8(32'hbb517ee4),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9da970),
	.w1(32'h3acf23d4),
	.w2(32'h3c347f70),
	.w3(32'h3bdd3367),
	.w4(32'h3babd87c),
	.w5(32'h3c5af6f4),
	.w6(32'hbb4e7898),
	.w7(32'h3b82dac6),
	.w8(32'hbb9583ba),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38fe99bf),
	.w1(32'hbbeb1ddb),
	.w2(32'hbba7a206),
	.w3(32'h3b196527),
	.w4(32'hbb364095),
	.w5(32'hbb703ef9),
	.w6(32'hbc167b46),
	.w7(32'hbbd46752),
	.w8(32'hbbbdf63b),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba77a020),
	.w1(32'hbab32bcc),
	.w2(32'hbb3425f7),
	.w3(32'h3b0efcf8),
	.w4(32'hbba86101),
	.w5(32'hbc06780a),
	.w6(32'h3b968777),
	.w7(32'hbbb02e82),
	.w8(32'hbc666684),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa45013),
	.w1(32'h3c274404),
	.w2(32'hb99a1e84),
	.w3(32'h3b8def20),
	.w4(32'h3c880f3d),
	.w5(32'h3c1c066f),
	.w6(32'h3b875a14),
	.w7(32'h3c91e731),
	.w8(32'h3c34d297),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc0db82),
	.w1(32'h3b22f70c),
	.w2(32'hbb931417),
	.w3(32'hbb85b5cc),
	.w4(32'h392c0e8e),
	.w5(32'hbc07e8ea),
	.w6(32'hbb07fd1f),
	.w7(32'h3bd013fc),
	.w8(32'hbb8aa156),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba03ab2),
	.w1(32'h3a00813e),
	.w2(32'hbb391b48),
	.w3(32'hbb5ae097),
	.w4(32'h3b0b8b06),
	.w5(32'h39a43d5c),
	.w6(32'hbb79e99d),
	.w7(32'hbab06927),
	.w8(32'hbb8c51f0),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9d920d),
	.w1(32'h3bee5e7f),
	.w2(32'h3b93121b),
	.w3(32'h3b6d9718),
	.w4(32'h3c302ac7),
	.w5(32'h3bd57b78),
	.w6(32'hbaa49304),
	.w7(32'h3b49e287),
	.w8(32'h3c1fcdfc),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba220d8f),
	.w1(32'hbc2dc9ea),
	.w2(32'hba5a3d2c),
	.w3(32'h39bc14f0),
	.w4(32'hbc00d106),
	.w5(32'hbb170d0b),
	.w6(32'h3b8086a5),
	.w7(32'hbbcd7df9),
	.w8(32'h3a83d3d6),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb969ca6),
	.w1(32'hba2cec6d),
	.w2(32'hbb24f84e),
	.w3(32'h3ba4fdbd),
	.w4(32'hbbe1ba32),
	.w5(32'hbb034e60),
	.w6(32'h3b1c455a),
	.w7(32'hbb569446),
	.w8(32'hbb67b60e),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3431ea),
	.w1(32'hb9ddead1),
	.w2(32'h3a6c021c),
	.w3(32'hbb0eae3e),
	.w4(32'hbbdb12a4),
	.w5(32'hbb8ee7f3),
	.w6(32'hbb856f1f),
	.w7(32'hbbf3abcb),
	.w8(32'hbba6765d),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baa26b9),
	.w1(32'hbac0ce32),
	.w2(32'hba96ba84),
	.w3(32'h3ba0fe83),
	.w4(32'h3a79d13d),
	.w5(32'hbb93f415),
	.w6(32'h3bd104c6),
	.w7(32'h391a5735),
	.w8(32'hbc386a95),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc857713),
	.w1(32'hbc08ef4f),
	.w2(32'hbc8ce702),
	.w3(32'hbc58be78),
	.w4(32'hbc06bcea),
	.w5(32'hbc0a8589),
	.w6(32'hbc32a965),
	.w7(32'hb9a04e7b),
	.w8(32'hbb17c4af),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5e7901),
	.w1(32'hbbc60d98),
	.w2(32'hbb7482c7),
	.w3(32'hbc63528a),
	.w4(32'hbc157575),
	.w5(32'hbc3fd6ec),
	.w6(32'hbc28f2ae),
	.w7(32'hbb8cb3ad),
	.w8(32'hbb827648),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbcbd1c),
	.w1(32'hbae9e84f),
	.w2(32'hbb020b66),
	.w3(32'h3b2c61b1),
	.w4(32'hbb593b86),
	.w5(32'hbab69cb4),
	.w6(32'h3a4fd745),
	.w7(32'hbb009693),
	.w8(32'h398c77cf),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b202a7c),
	.w1(32'h3b0ca04a),
	.w2(32'hbb439024),
	.w3(32'h3baf3218),
	.w4(32'h3b8f644e),
	.w5(32'hba4416c7),
	.w6(32'h3bf14d1c),
	.w7(32'h3b44dcc7),
	.w8(32'hbb714173),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafa282d),
	.w1(32'hba8c26ab),
	.w2(32'hb9629cab),
	.w3(32'hbb13f2ab),
	.w4(32'hbc101a3c),
	.w5(32'h3bc86616),
	.w6(32'hbb6fd32b),
	.w7(32'hbbf1cb67),
	.w8(32'hbbbf18a9),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9fc357),
	.w1(32'h3bd902cc),
	.w2(32'hb95e1d46),
	.w3(32'hbbaacc9b),
	.w4(32'h3a479a9d),
	.w5(32'h3c24a3aa),
	.w6(32'hbb07036f),
	.w7(32'h3aed446f),
	.w8(32'hbac4bb79),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c80741d),
	.w1(32'h3c4a6e83),
	.w2(32'h3c77dc87),
	.w3(32'h3c875504),
	.w4(32'h3c9aa232),
	.w5(32'h3bef127e),
	.w6(32'h3c8fbdee),
	.w7(32'h3c8c52e6),
	.w8(32'h3c582f01),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1b158d),
	.w1(32'h3b105ba5),
	.w2(32'h395011f6),
	.w3(32'h3bbba671),
	.w4(32'h3ad0488b),
	.w5(32'h3b01c0c1),
	.w6(32'h3c1d3cf1),
	.w7(32'h3ac737b1),
	.w8(32'h3b328356),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1bdb33),
	.w1(32'h3c2bcca5),
	.w2(32'h3b61c621),
	.w3(32'h3c08fd8a),
	.w4(32'h3bf66ed5),
	.w5(32'h3b25df16),
	.w6(32'h3c38ede9),
	.w7(32'h3c2291f2),
	.w8(32'h3b932e93),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abe02cd),
	.w1(32'h3b80d72b),
	.w2(32'h3bf4976a),
	.w3(32'hbb69d4b6),
	.w4(32'hbb29ecb5),
	.w5(32'h3b936699),
	.w6(32'hbb0ad548),
	.w7(32'hba5832bd),
	.w8(32'hba511e2d),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cafaf90),
	.w1(32'hbb9b7ec0),
	.w2(32'h3ae370bc),
	.w3(32'h3cc5bfed),
	.w4(32'h3b74c150),
	.w5(32'h3c469d93),
	.w6(32'h3c7c67e4),
	.w7(32'h3b86744f),
	.w8(32'h3bc11797),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb329798),
	.w1(32'hbb9a24fa),
	.w2(32'h3bb2972b),
	.w3(32'hbb84ffba),
	.w4(32'hbc0acf9d),
	.w5(32'hbb235e7d),
	.w6(32'hbaebfc06),
	.w7(32'hbabb6e94),
	.w8(32'hb92f84cc),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d8a4db),
	.w1(32'h3b231867),
	.w2(32'h3b993716),
	.w3(32'h3ae925f1),
	.w4(32'hba7d84af),
	.w5(32'h3994d399),
	.w6(32'hbacf51bf),
	.w7(32'hbb587f53),
	.w8(32'hbb07b6af),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1c84a5),
	.w1(32'hb9e4a8cc),
	.w2(32'hbb3fa3b6),
	.w3(32'h3b309f12),
	.w4(32'hb9d9d8ac),
	.w5(32'hbb01ecd1),
	.w6(32'h3b195e44),
	.w7(32'hb91b25b0),
	.w8(32'h3af6afa2),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c248275),
	.w1(32'h3baa909e),
	.w2(32'h3b833099),
	.w3(32'h3c1dfd87),
	.w4(32'h3be25a23),
	.w5(32'h3c9027f2),
	.w6(32'h3c21a027),
	.w7(32'h3c830881),
	.w8(32'h3c8aafc6),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc0ac4b),
	.w1(32'hba8228a3),
	.w2(32'h3bc9b782),
	.w3(32'hbbbdc408),
	.w4(32'hbc1588e3),
	.w5(32'h395cae64),
	.w6(32'hbbd48a60),
	.w7(32'hbb9e3105),
	.w8(32'hbb0bfb15),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfe7563),
	.w1(32'h3bd2d85b),
	.w2(32'h3c7c17f8),
	.w3(32'h3c57c8d8),
	.w4(32'hb9014de4),
	.w5(32'h3c4475c9),
	.w6(32'h3ac4bba6),
	.w7(32'hbad5001d),
	.w8(32'h3bb3e224),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba213fcc),
	.w1(32'hbb31781c),
	.w2(32'hbb7d7e66),
	.w3(32'h3b87cac4),
	.w4(32'hba99e86b),
	.w5(32'hbaba94bb),
	.w6(32'h3b818269),
	.w7(32'h3a8d0b1d),
	.w8(32'h3b16fe8f),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba3ecf7),
	.w1(32'h3bc1166b),
	.w2(32'h3b55972a),
	.w3(32'h3c044b3a),
	.w4(32'h3b7ae79e),
	.w5(32'h3c19ed7b),
	.w6(32'h3c226e81),
	.w7(32'h3bf941b3),
	.w8(32'h3bd6b43f),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f1527d),
	.w1(32'hbb8a6029),
	.w2(32'hbabd0aaa),
	.w3(32'h3b83aeb6),
	.w4(32'hb9226335),
	.w5(32'h3bbe3350),
	.w6(32'h3ba955a4),
	.w7(32'hbae714dd),
	.w8(32'h3b069c77),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac134dc),
	.w1(32'h3ba8548d),
	.w2(32'h3b5487c9),
	.w3(32'hbb913b24),
	.w4(32'hba803b90),
	.w5(32'h3c92b6d1),
	.w6(32'hbab21644),
	.w7(32'hbc15e743),
	.w8(32'h3c3bcc8a),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3086b9),
	.w1(32'hbb9ef38e),
	.w2(32'hbbd630fd),
	.w3(32'hb9c92c5e),
	.w4(32'hbb2da92d),
	.w5(32'hbb8d2b56),
	.w6(32'h3b161429),
	.w7(32'hbb0cf873),
	.w8(32'hbc04cc45),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0d6964),
	.w1(32'hbba5a400),
	.w2(32'hbadaaebe),
	.w3(32'h3b7fd93b),
	.w4(32'hbb38bb66),
	.w5(32'h3b56c597),
	.w6(32'h3885b7e7),
	.w7(32'hbbbac2ac),
	.w8(32'hbb06e575),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4a4396),
	.w1(32'hbb424b5e),
	.w2(32'h3c6e1741),
	.w3(32'h3c473a11),
	.w4(32'h3a152505),
	.w5(32'h3c01493f),
	.w6(32'h3b16591d),
	.w7(32'h3bbe15f7),
	.w8(32'h3b7e5c71),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c67e21c),
	.w1(32'h39a408c7),
	.w2(32'h3bc388ac),
	.w3(32'h3ba91899),
	.w4(32'h3b2e637c),
	.w5(32'h3ba4c051),
	.w6(32'h3a8a2fd4),
	.w7(32'h3a9727bf),
	.w8(32'h3c0d8c48),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8a3a95),
	.w1(32'h3b8087c5),
	.w2(32'hbabc3ad2),
	.w3(32'hbadad929),
	.w4(32'h3a8874a2),
	.w5(32'hbb17ce05),
	.w6(32'hba503a2c),
	.w7(32'h3aacf497),
	.w8(32'hbc03916a),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbace5ec0),
	.w1(32'h3b2f912a),
	.w2(32'h3a32d459),
	.w3(32'hbba14b56),
	.w4(32'h3bd86ffe),
	.w5(32'hb9a47b2d),
	.w6(32'hbb1e8c75),
	.w7(32'h3b45c781),
	.w8(32'h3b64001c),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38819564),
	.w1(32'h3c09935e),
	.w2(32'h3b99e1cf),
	.w3(32'hba4fd9aa),
	.w4(32'h3c24bf64),
	.w5(32'h3b49c768),
	.w6(32'h3b670d25),
	.w7(32'h3c11dd52),
	.w8(32'h3bc02a6c),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b43d1fb),
	.w1(32'hbbd27b4e),
	.w2(32'h3b11ca54),
	.w3(32'h3ac6afa2),
	.w4(32'hbc207292),
	.w5(32'hbad501ff),
	.w6(32'h3b93451c),
	.w7(32'hbb8a3110),
	.w8(32'hbbbd4f53),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98425b5),
	.w1(32'hbbd1e1be),
	.w2(32'h3b841d8e),
	.w3(32'h39dba76a),
	.w4(32'hbb93d017),
	.w5(32'h3bb50db4),
	.w6(32'hbc1e0396),
	.w7(32'hbc2fb8ee),
	.w8(32'hbb00972f),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b914570),
	.w1(32'h3c29a2f1),
	.w2(32'h3c398174),
	.w3(32'hba919c0c),
	.w4(32'h3b21ecda),
	.w5(32'hb8b38a38),
	.w6(32'hbac1aa80),
	.w7(32'h3c094368),
	.w8(32'h3c1b48ab),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afe8841),
	.w1(32'h3a7ce98f),
	.w2(32'h3b30fc22),
	.w3(32'hbb987c6a),
	.w4(32'h3ad41e41),
	.w5(32'h3b74675f),
	.w6(32'hbb5f0668),
	.w7(32'hbad6dbb9),
	.w8(32'h3a708ee7),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbddc676),
	.w1(32'hbb4c87fd),
	.w2(32'hbc4049df),
	.w3(32'hbb6c2788),
	.w4(32'hbc110cd0),
	.w5(32'hbc4f6b45),
	.w6(32'hbb5bd4ef),
	.w7(32'hbc349332),
	.w8(32'h3b1dcebe),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7790cf),
	.w1(32'h3bdb442d),
	.w2(32'h3b70f844),
	.w3(32'hbbf54da5),
	.w4(32'hbc682c11),
	.w5(32'hbc373c9d),
	.w6(32'hbbcfcd2a),
	.w7(32'hbae7970f),
	.w8(32'hbc125a57),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9d97a3),
	.w1(32'h3b13be8d),
	.w2(32'h3c786db1),
	.w3(32'hbc01ab6d),
	.w4(32'h3c0bc91d),
	.w5(32'h3c3f9953),
	.w6(32'hba355a22),
	.w7(32'h3ae019e3),
	.w8(32'h3aae3e79),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b2c588),
	.w1(32'h395633d7),
	.w2(32'hbc78180f),
	.w3(32'h3c186035),
	.w4(32'h3ae4f213),
	.w5(32'hbb0ccd58),
	.w6(32'hba8175a9),
	.w7(32'h3b850b14),
	.w8(32'h3b95a573),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc65e253),
	.w1(32'h3b17db8d),
	.w2(32'h3b0453ff),
	.w3(32'hbb193c05),
	.w4(32'h3c3e7c3f),
	.w5(32'h3c290b99),
	.w6(32'hbb43aeda),
	.w7(32'h3bdb989f),
	.w8(32'h3be40be5),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b30b9d1),
	.w1(32'h3b25f98e),
	.w2(32'hbb93957a),
	.w3(32'h3b0f0613),
	.w4(32'h3c2ed4e4),
	.w5(32'h3d515f77),
	.w6(32'h39e22246),
	.w7(32'hbae3b37d),
	.w8(32'hbb18ac8b),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be5ac15),
	.w1(32'h3c19c072),
	.w2(32'h3c558dd8),
	.w3(32'h3c9c0e1d),
	.w4(32'h3beaa948),
	.w5(32'h3cbbc342),
	.w6(32'h3c1575cc),
	.w7(32'hbc127704),
	.w8(32'h3a82c671),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc20174),
	.w1(32'h3b34ea4a),
	.w2(32'h3ba7294c),
	.w3(32'h3c16e885),
	.w4(32'hbaa448d4),
	.w5(32'hb9876f0c),
	.w6(32'h3bf997f4),
	.w7(32'hbbd8a1ed),
	.w8(32'hbc5f97e5),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c829dc1),
	.w1(32'h3c3cb355),
	.w2(32'h3c8110b6),
	.w3(32'h3c16797f),
	.w4(32'h3c945c60),
	.w5(32'h3c9bbe58),
	.w6(32'h3afb73ad),
	.w7(32'h3bebc493),
	.w8(32'h3c1ba4ec),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfa3f8f),
	.w1(32'hbb99378c),
	.w2(32'h3ba5d696),
	.w3(32'h3c8d9f75),
	.w4(32'hba172064),
	.w5(32'h3beefbcb),
	.w6(32'h3c245741),
	.w7(32'hbc2b5421),
	.w8(32'hbab6dfa2),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3d0ef3),
	.w1(32'hbb80fe59),
	.w2(32'hbc0237e1),
	.w3(32'h3b9d7e83),
	.w4(32'hbb856d94),
	.w5(32'hbba0a76e),
	.w6(32'hbb1c065a),
	.w7(32'h3c019be5),
	.w8(32'hbc94a81f),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca71e6f),
	.w1(32'h3baf8375),
	.w2(32'h3c017097),
	.w3(32'h3ad9cbe2),
	.w4(32'hbc074162),
	.w5(32'hbc85e541),
	.w6(32'hbb52f142),
	.w7(32'h3bed0f43),
	.w8(32'h3bc69fa5),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8f4fcf),
	.w1(32'h3b1c8d39),
	.w2(32'h3c0812b7),
	.w3(32'h3b80f1bd),
	.w4(32'h3ab9070c),
	.w5(32'h3b61f6d8),
	.w6(32'h3c4c3da8),
	.w7(32'h3b0b64b8),
	.w8(32'hba869ca8),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf02f99),
	.w1(32'h3af7d820),
	.w2(32'h3b928047),
	.w3(32'h3c12561a),
	.w4(32'h3b51cab7),
	.w5(32'h3b95efdd),
	.w6(32'h3944969e),
	.w7(32'hbb0ff351),
	.w8(32'hbb355b61),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd696b8),
	.w1(32'hba9c78f1),
	.w2(32'hbc2bbcc1),
	.w3(32'h3c046f32),
	.w4(32'hbb4f3bbf),
	.w5(32'hbba604a2),
	.w6(32'h3b8eb00a),
	.w7(32'h38b28074),
	.w8(32'hbbcbda3f),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0a2b97),
	.w1(32'h3b8896ce),
	.w2(32'h3cad1468),
	.w3(32'h3a7e1c93),
	.w4(32'h3a57b8d2),
	.w5(32'h3c08cadd),
	.w6(32'hbbf999b5),
	.w7(32'hba3fbf02),
	.w8(32'h3b8b0078),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b63d4b7),
	.w1(32'hbc63339d),
	.w2(32'hbc03e504),
	.w3(32'h3c47abcb),
	.w4(32'hbbbc0002),
	.w5(32'hbc3cae9d),
	.w6(32'h3bcdcf59),
	.w7(32'h3a326a1e),
	.w8(32'hb8e2dd89),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb99b838),
	.w1(32'hbb38992d),
	.w2(32'hbaf7c545),
	.w3(32'hbc07b09f),
	.w4(32'hbc395879),
	.w5(32'hbba16197),
	.w6(32'h3b90fb1e),
	.w7(32'h3c0cd6ee),
	.w8(32'h39967f22),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c30556b),
	.w1(32'hbb3eaa0b),
	.w2(32'hbba759f8),
	.w3(32'h3ada835f),
	.w4(32'hbabbe98a),
	.w5(32'h3c75a927),
	.w6(32'h3a85142e),
	.w7(32'hbc04164f),
	.w8(32'hb627d294),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb06323e),
	.w1(32'h3b41bc68),
	.w2(32'h3bb0aa30),
	.w3(32'h3bb53506),
	.w4(32'hbb882cd7),
	.w5(32'hbb9cf364),
	.w6(32'h3be5d688),
	.w7(32'hbbbd3f2c),
	.w8(32'hbc028bcf),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b14e3a0),
	.w1(32'h3c1cae44),
	.w2(32'h3b41659f),
	.w3(32'h3a32c1fc),
	.w4(32'h3c6b94e2),
	.w5(32'hba8f7fec),
	.w6(32'hbbcdead1),
	.w7(32'h3c18c9f4),
	.w8(32'h3c0521ab),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1aa35a),
	.w1(32'hbbe18d2e),
	.w2(32'h39907a9e),
	.w3(32'hbc69b3e6),
	.w4(32'hbbe6a53d),
	.w5(32'hbc6be9c4),
	.w6(32'hbc476f3f),
	.w7(32'hbb98df66),
	.w8(32'hbbfbee0d),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdeee0f),
	.w1(32'hbc58d7ee),
	.w2(32'hbc63314d),
	.w3(32'h3c01ae93),
	.w4(32'hbc49f8d6),
	.w5(32'hbc00fd2d),
	.w6(32'h3b479c26),
	.w7(32'h3aee5616),
	.w8(32'hbb271fa8),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9f42f4),
	.w1(32'hbc4f2433),
	.w2(32'hbc7cf73e),
	.w3(32'hbc8cd5a8),
	.w4(32'hbad9933c),
	.w5(32'h3a281bb7),
	.w6(32'h3b1e58aa),
	.w7(32'hbbb2702a),
	.w8(32'hbc08ecce),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb698efe),
	.w1(32'hbb7b6f89),
	.w2(32'hbb307999),
	.w3(32'h3b155c20),
	.w4(32'hbc012ae1),
	.w5(32'hbb217ff9),
	.w6(32'hbb55873f),
	.w7(32'hbbc29f62),
	.w8(32'hbb421d64),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7cad9e),
	.w1(32'h3b88dd27),
	.w2(32'h3afaf725),
	.w3(32'hbc1d2e2b),
	.w4(32'hbc936eef),
	.w5(32'hbc00aff3),
	.w6(32'hbbadba4a),
	.w7(32'hbb8b141c),
	.w8(32'hbc926941),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c25006a),
	.w1(32'hbc0ce5ed),
	.w2(32'hbc67019a),
	.w3(32'hbc802b86),
	.w4(32'h3ae76f6d),
	.w5(32'hbb3c971a),
	.w6(32'hbc012514),
	.w7(32'h3a1b0f08),
	.w8(32'hbc07590a),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5046b3),
	.w1(32'hbb5910a4),
	.w2(32'hbbc418b7),
	.w3(32'h3aac49ca),
	.w4(32'hbbfadbbf),
	.w5(32'hbb2731ea),
	.w6(32'hbc84074d),
	.w7(32'hbbab4e97),
	.w8(32'hbb4720c2),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8f9121),
	.w1(32'h3c4932f4),
	.w2(32'h3b4084f9),
	.w3(32'hbac4e2f0),
	.w4(32'h3b8190cd),
	.w5(32'hb996a55b),
	.w6(32'h399a6ab1),
	.w7(32'hbc07cde9),
	.w8(32'h3b84e2e6),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdec04a),
	.w1(32'hbc30c4cb),
	.w2(32'hbbb7badb),
	.w3(32'hbc67d162),
	.w4(32'hbb47adb2),
	.w5(32'hbc3ac82b),
	.w6(32'hbc9829c5),
	.w7(32'hbc110923),
	.w8(32'hbb231e7c),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb41b002),
	.w1(32'h3b1dd652),
	.w2(32'hbbe71c99),
	.w3(32'hbbc9a4f8),
	.w4(32'h3ce0e687),
	.w5(32'h3d085c28),
	.w6(32'hbbd8c66a),
	.w7(32'h3c30e9ae),
	.w8(32'h3c7b657d),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb40a68),
	.w1(32'hbb342e92),
	.w2(32'hbc66ba0b),
	.w3(32'h3c7bc624),
	.w4(32'hbc3a8671),
	.w5(32'hbc762332),
	.w6(32'h3bcbf8b8),
	.w7(32'hbc4f350f),
	.w8(32'hbca4a292),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9b9bd7),
	.w1(32'h3b32ec39),
	.w2(32'hbb49e934),
	.w3(32'h3be59a6b),
	.w4(32'h3bb9f780),
	.w5(32'h3c5069ad),
	.w6(32'h3c26212d),
	.w7(32'hbb24dad8),
	.w8(32'hba98a941),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc59fe3a),
	.w1(32'hbb4e9713),
	.w2(32'h3b9e0fa6),
	.w3(32'h3af85b1d),
	.w4(32'h3c5a63b6),
	.w5(32'h3c1dda87),
	.w6(32'hba10c6d6),
	.w7(32'hbbdbfecc),
	.w8(32'hbbfae7ec),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39aecd8d),
	.w1(32'hbb363060),
	.w2(32'h3af3c090),
	.w3(32'h3ba8f547),
	.w4(32'hbbb8669e),
	.w5(32'h3a946f57),
	.w6(32'hbbc1a209),
	.w7(32'hbc12bb0f),
	.w8(32'hbb99215f),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c051274),
	.w1(32'h3b0775c9),
	.w2(32'h3a6f64df),
	.w3(32'h3baa660e),
	.w4(32'hbc33180d),
	.w5(32'hbb817f9a),
	.w6(32'hbb7e6e48),
	.w7(32'hbba0aeae),
	.w8(32'hbc162461),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aebd679),
	.w1(32'hbc291941),
	.w2(32'hbc057309),
	.w3(32'hbc6c8187),
	.w4(32'hbba1f89b),
	.w5(32'hbb8450aa),
	.w6(32'hbb5133b5),
	.w7(32'hb9ea234a),
	.w8(32'h3bacc108),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3943da45),
	.w1(32'h3bc9a848),
	.w2(32'h3b3651ae),
	.w3(32'hb9f1096f),
	.w4(32'h3b79a569),
	.w5(32'h3aa653f7),
	.w6(32'h3c1176b2),
	.w7(32'hbb167ed9),
	.w8(32'hbb5e2e6b),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc196ce),
	.w1(32'h3bd83496),
	.w2(32'hba23d573),
	.w3(32'hba101412),
	.w4(32'h3c80c867),
	.w5(32'h3bc66e82),
	.w6(32'h3b90dc59),
	.w7(32'h3c1c05b1),
	.w8(32'h3bac01ad),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fc4986),
	.w1(32'h3ac05993),
	.w2(32'h3b4158fb),
	.w3(32'h3c690fbd),
	.w4(32'h3c328912),
	.w5(32'h3c4a2d01),
	.w6(32'h3c9057c5),
	.w7(32'h3b458165),
	.w8(32'h3c3ced25),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b910e59),
	.w1(32'hbb395d86),
	.w2(32'hbc104f67),
	.w3(32'h3c73ff8b),
	.w4(32'hbb413d8c),
	.w5(32'h3c16b2ae),
	.w6(32'h3c243604),
	.w7(32'h3bf54e17),
	.w8(32'hbc1aac77),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc8894a),
	.w1(32'hbc0bcef7),
	.w2(32'hbb31a32a),
	.w3(32'hbc756713),
	.w4(32'h3b54ff7d),
	.w5(32'h3b10b8c0),
	.w6(32'hbbdf8b7b),
	.w7(32'h3bf22d43),
	.w8(32'h3a664bdc),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad42359),
	.w1(32'h3bbbd28b),
	.w2(32'h3ada4e98),
	.w3(32'hbad66c3f),
	.w4(32'h3c121a6f),
	.w5(32'h3a958401),
	.w6(32'hbbe56dc2),
	.w7(32'h3c94db57),
	.w8(32'h3c5a3da3),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b90b324),
	.w1(32'hba81389e),
	.w2(32'hbb223067),
	.w3(32'hbacb64fd),
	.w4(32'hbb1d6d48),
	.w5(32'h3b82bf3d),
	.w6(32'h3c01c7bf),
	.w7(32'h3b2c50a7),
	.w8(32'h3bcf041e),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2f1f88),
	.w1(32'h3c2fb9bd),
	.w2(32'h3ca054ee),
	.w3(32'h3c412256),
	.w4(32'h3c1fd22d),
	.w5(32'h3c0f4c74),
	.w6(32'h3c722465),
	.w7(32'hbac8236c),
	.w8(32'hbaed84e6),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b347504),
	.w1(32'hbc2d442c),
	.w2(32'hbb55b512),
	.w3(32'h3a9b83e2),
	.w4(32'h39f70c0a),
	.w5(32'hba9a02d7),
	.w6(32'h39c0c5b1),
	.w7(32'h3bc8fbed),
	.w8(32'h3bf4b26c),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb57420c),
	.w1(32'hba983693),
	.w2(32'hba8b37a7),
	.w3(32'hbb47a426),
	.w4(32'hbb669f77),
	.w5(32'hbb116e9f),
	.w6(32'h3bbd4283),
	.w7(32'hbbd1812a),
	.w8(32'hbbade137),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b84df8a),
	.w1(32'h39e4e7f4),
	.w2(32'h3a96fcfd),
	.w3(32'h3becfbd1),
	.w4(32'hbc06c892),
	.w5(32'hbb8058a5),
	.w6(32'h3c2edf43),
	.w7(32'hbc09a1bf),
	.w8(32'hbc0b1e51),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7ba9a3),
	.w1(32'h3b2cfad9),
	.w2(32'hbb3e7a4d),
	.w3(32'h3b00b439),
	.w4(32'hbb8460e6),
	.w5(32'hbc769aa3),
	.w6(32'hbba77103),
	.w7(32'hbbe97492),
	.w8(32'hbb1ab905),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bab7837),
	.w1(32'h3b2df7fb),
	.w2(32'h3b3ff0bf),
	.w3(32'hbb505843),
	.w4(32'h3bcce70e),
	.w5(32'h3c2d01cb),
	.w6(32'hba0074e5),
	.w7(32'hbbc034dd),
	.w8(32'hbb50a43f),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b01a9c2),
	.w1(32'hbb60a395),
	.w2(32'hbb689de6),
	.w3(32'h3c5f54a9),
	.w4(32'h3ae75033),
	.w5(32'hbbd52a34),
	.w6(32'h3ba472f6),
	.w7(32'h3b8552a2),
	.w8(32'hbb040292),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc10f7c1),
	.w1(32'hbbbf632a),
	.w2(32'hbb545aad),
	.w3(32'hbc1632e8),
	.w4(32'hbb89cc72),
	.w5(32'hbbf67910),
	.w6(32'hbbf2a3e2),
	.w7(32'hbbd6ce28),
	.w8(32'hbc277316),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2ce1c5),
	.w1(32'hbc56099f),
	.w2(32'hbc0d85f3),
	.w3(32'h3ae3099f),
	.w4(32'hbbed8159),
	.w5(32'hbc1f2713),
	.w6(32'hbb90b3ec),
	.w7(32'h3b43d158),
	.w8(32'h3c826982),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf2a4d9),
	.w1(32'h3bdaf95a),
	.w2(32'h3b1f6f8b),
	.w3(32'h3c4ad5c9),
	.w4(32'hb8f3da25),
	.w5(32'h3b7e0979),
	.w6(32'h3c083e8b),
	.w7(32'h3bb904ef),
	.w8(32'h3ba05496),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bad0933),
	.w1(32'h3a22762f),
	.w2(32'h3beb5188),
	.w3(32'h3891a529),
	.w4(32'h3bbad02d),
	.w5(32'h3bc52069),
	.w6(32'h3a9ca22d),
	.w7(32'hbb3df716),
	.w8(32'h3b95a5d0),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb35267e),
	.w1(32'h3b5de07d),
	.w2(32'h3c721ebf),
	.w3(32'h3bbe465f),
	.w4(32'h3bd6b245),
	.w5(32'h3c3845b5),
	.w6(32'h3c05f37b),
	.w7(32'hbbcd625c),
	.w8(32'hba74f965),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb732f61),
	.w1(32'h3c0d43eb),
	.w2(32'h3b8cc646),
	.w3(32'h3c2add7c),
	.w4(32'hb99fae97),
	.w5(32'h3b86befe),
	.w6(32'h396dcec0),
	.w7(32'hba732bf2),
	.w8(32'hbb9eb946),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a99a327),
	.w1(32'hbc0bfd4f),
	.w2(32'h3c27622b),
	.w3(32'hba0b27a8),
	.w4(32'hbc2f19d5),
	.w5(32'h3bfe283b),
	.w6(32'h3b0cf7c5),
	.w7(32'h3c17d6e1),
	.w8(32'h3bf81287),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2baacc),
	.w1(32'hbb33dc1b),
	.w2(32'hbb845f52),
	.w3(32'hbafc2688),
	.w4(32'hbbd84033),
	.w5(32'h3ac18517),
	.w6(32'h3a461766),
	.w7(32'hbb33690c),
	.w8(32'hbb85c0a9),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb946c60),
	.w1(32'h3bea64a2),
	.w2(32'h3c33a90f),
	.w3(32'hbad68190),
	.w4(32'h3afc55fc),
	.w5(32'h3c3c4973),
	.w6(32'hb9c0e3d2),
	.w7(32'h3c797f4f),
	.w8(32'h3bc79acc),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd8fef0),
	.w1(32'h3ba544ff),
	.w2(32'h3bd51fba),
	.w3(32'h380553c7),
	.w4(32'h3b28e778),
	.w5(32'h3bf61135),
	.w6(32'h3a9a8b37),
	.w7(32'hbbd65b6f),
	.w8(32'hbbcbd709),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9870879),
	.w1(32'h3acbeea1),
	.w2(32'hbb6355c2),
	.w3(32'h3a83968c),
	.w4(32'h390297e3),
	.w5(32'h3c670b83),
	.w6(32'h3b58fc3c),
	.w7(32'hbb38528a),
	.w8(32'h3a5e92fe),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba95a3b6),
	.w1(32'hbbcbea69),
	.w2(32'hbc2d5077),
	.w3(32'hbbda63a6),
	.w4(32'hbbc999df),
	.w5(32'hbb38fd6c),
	.w6(32'hbb4d578f),
	.w7(32'h3bd649d9),
	.w8(32'h3b95d5be),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b97383a),
	.w1(32'h3bfff19e),
	.w2(32'h3bdc3e99),
	.w3(32'h3b949364),
	.w4(32'h3c2690b0),
	.w5(32'h3bf29567),
	.w6(32'h3b8f14ce),
	.w7(32'h3b363fba),
	.w8(32'h3c1afe9d),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb42324),
	.w1(32'h3b589588),
	.w2(32'h3c3f9159),
	.w3(32'h3b4176eb),
	.w4(32'h3c38eb94),
	.w5(32'h3c180038),
	.w6(32'h3bf31845),
	.w7(32'hbb564f1c),
	.w8(32'h3a89fefa),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb6627a),
	.w1(32'h3c162437),
	.w2(32'h3c7e848a),
	.w3(32'hbb217f1c),
	.w4(32'h3c32e523),
	.w5(32'h3c3fe572),
	.w6(32'h3b7f7443),
	.w7(32'hbb15d8c4),
	.w8(32'h3ba1a00a),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd3e534),
	.w1(32'hbb4dabb9),
	.w2(32'hbc11142c),
	.w3(32'h3c234fc8),
	.w4(32'hbabdcd14),
	.w5(32'hbc3ee74f),
	.w6(32'hbae8a3ef),
	.w7(32'hba36c2f3),
	.w8(32'hbb5c4f72),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be7cff7),
	.w1(32'h3ab337d6),
	.w2(32'hbad7f678),
	.w3(32'hbbcd679e),
	.w4(32'hbb7173a3),
	.w5(32'hbb504d36),
	.w6(32'hbbcf2e81),
	.w7(32'h3b064197),
	.w8(32'h3bc72a43),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f9f4be),
	.w1(32'h3bbc14a2),
	.w2(32'h3c1ef032),
	.w3(32'hbab47b1d),
	.w4(32'h3c5e4a77),
	.w5(32'h3c8a04cd),
	.w6(32'h3b8754d4),
	.w7(32'hbac11fb0),
	.w8(32'h3bbd59c6),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba9c8fe),
	.w1(32'hbbc6c524),
	.w2(32'hbb2da785),
	.w3(32'h3b63679e),
	.w4(32'h3ae4b755),
	.w5(32'h3c5d2240),
	.w6(32'h3bbc385a),
	.w7(32'hbb96391a),
	.w8(32'hbb777270),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5e62d0),
	.w1(32'h39c605c7),
	.w2(32'h3b94f102),
	.w3(32'h3c277bc8),
	.w4(32'h3983dc2e),
	.w5(32'hbb1b6ca5),
	.w6(32'h38cae01a),
	.w7(32'hbc22da1b),
	.w8(32'hbb1bf723),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa1b9e9),
	.w1(32'hbbbc7598),
	.w2(32'h3b508078),
	.w3(32'h3bde216f),
	.w4(32'hbc407408),
	.w5(32'hbbf63612),
	.w6(32'hba18f9d0),
	.w7(32'hbbe2dd8c),
	.w8(32'hbb07d4d6),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc94df7),
	.w1(32'h3ba541fc),
	.w2(32'hbbbe69f6),
	.w3(32'hbaada56d),
	.w4(32'h3c190292),
	.w5(32'h3c5b5dcd),
	.w6(32'h390c0bf2),
	.w7(32'h3bddd406),
	.w8(32'h3c0f1602),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb84fad6),
	.w1(32'h3c0535b2),
	.w2(32'h3c99156e),
	.w3(32'h3a990c69),
	.w4(32'hbb1869fd),
	.w5(32'h3c370976),
	.w6(32'h3b07c810),
	.w7(32'h3ba00943),
	.w8(32'h3bc96050),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb237430),
	.w1(32'h3b86edde),
	.w2(32'h3c30fab6),
	.w3(32'h3c383e17),
	.w4(32'h3b8f7aa4),
	.w5(32'hbbb462bc),
	.w6(32'h3b6d9f8a),
	.w7(32'hbb0affad),
	.w8(32'h397c867a),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb559617),
	.w1(32'h3c9ec6e3),
	.w2(32'h3d031f9c),
	.w3(32'h3b5c6237),
	.w4(32'h3c21e83d),
	.w5(32'h3a434495),
	.w6(32'hba47072b),
	.w7(32'hbb935261),
	.w8(32'h3a1a7be3),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c87fdaf),
	.w1(32'h3c3facae),
	.w2(32'h3bf09c41),
	.w3(32'h3c9aa144),
	.w4(32'h3be1f915),
	.w5(32'hbb8fafd7),
	.w6(32'h3a48a382),
	.w7(32'hbbf77fe5),
	.w8(32'hbc5afef9),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9e170e),
	.w1(32'h3be9f2d3),
	.w2(32'h3c6203e3),
	.w3(32'hbc228f11),
	.w4(32'hbb721a56),
	.w5(32'hba30d7cc),
	.w6(32'hbc66c0d5),
	.w7(32'hbc1b9d70),
	.w8(32'hbb816e55),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ccbb581),
	.w1(32'h3bc4fc0e),
	.w2(32'h3cb65f7f),
	.w3(32'h3cd5ce67),
	.w4(32'h3c807052),
	.w5(32'h3ca0a07b),
	.w6(32'h3c4c0ad2),
	.w7(32'h3bbed24c),
	.w8(32'h3caee7f3),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb822b3),
	.w1(32'hbc082344),
	.w2(32'hbaadad88),
	.w3(32'h3cc6ac0f),
	.w4(32'hbb2ceec6),
	.w5(32'hbbf6ceed),
	.w6(32'h3c9fe0e4),
	.w7(32'hbb0a9131),
	.w8(32'hbb722307),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c04c0df),
	.w1(32'hbbf3ed7d),
	.w2(32'h3a20d0a1),
	.w3(32'h3b3476d2),
	.w4(32'hbb270fef),
	.w5(32'h3a470ea3),
	.w6(32'h3aff74f8),
	.w7(32'h3bda0a75),
	.w8(32'h3b5c7aed),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af9b7e2),
	.w1(32'hbbcdb271),
	.w2(32'hbadc65ee),
	.w3(32'hbb890f49),
	.w4(32'hbb666a3b),
	.w5(32'h3c0a3a9f),
	.w6(32'hbbd749eb),
	.w7(32'h3b247b1e),
	.w8(32'hbbd883f0),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c39e1a7),
	.w1(32'hbbc33bec),
	.w2(32'hbc7d8e83),
	.w3(32'h3c0ce201),
	.w4(32'hbb8c1e2e),
	.w5(32'hbc68a8f8),
	.w6(32'hbbbe7320),
	.w7(32'hba91325c),
	.w8(32'hbc1ae92c),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3304f8),
	.w1(32'hbc46ff3c),
	.w2(32'hbc863d5e),
	.w3(32'hbbf6e241),
	.w4(32'hbb9d8b36),
	.w5(32'hbc168724),
	.w6(32'h39ac0e49),
	.w7(32'h3c321753),
	.w8(32'h3c1293e9),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb750fac),
	.w1(32'hba7138c8),
	.w2(32'h3b8648e1),
	.w3(32'hbbc70144),
	.w4(32'hbaadd9fc),
	.w5(32'hbbe7aaf4),
	.w6(32'hbb827b3d),
	.w7(32'h3c016696),
	.w8(32'h3bab0b0a),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb23d5e9),
	.w1(32'hbbeda3fd),
	.w2(32'hbbbd7bcf),
	.w3(32'hbbd3eac9),
	.w4(32'hbc2cbd8a),
	.w5(32'hbc24ac60),
	.w6(32'h3ba05895),
	.w7(32'hbb1ece62),
	.w8(32'hba4cfff5),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8306c98),
	.w1(32'h3b4adb4c),
	.w2(32'hbb3b2f0a),
	.w3(32'hbb1c9493),
	.w4(32'hbb7a1cdf),
	.w5(32'hbb9a4604),
	.w6(32'h3b152890),
	.w7(32'hbb0e7763),
	.w8(32'h3b474f39),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2dd0d2),
	.w1(32'hba049a6d),
	.w2(32'h3c936ae0),
	.w3(32'hbb65b28f),
	.w4(32'h3c1a4831),
	.w5(32'h3bff506e),
	.w6(32'hbc03aea4),
	.w7(32'h3b7b012d),
	.w8(32'hbaaac287),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c63094d),
	.w1(32'h3ad9ecf8),
	.w2(32'hb9f57944),
	.w3(32'hbb8b55e7),
	.w4(32'h3bf4e7ca),
	.w5(32'h3b3c2ef8),
	.w6(32'hbbab68dc),
	.w7(32'hbb946474),
	.w8(32'hb9e4004b),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb74cdf4),
	.w1(32'h3c19eb88),
	.w2(32'h3cbe4e2f),
	.w3(32'h3b17cd00),
	.w4(32'h3c2d5412),
	.w5(32'hba863206),
	.w6(32'hbac961d2),
	.w7(32'hbbcd5718),
	.w8(32'hbb5b9112),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c99dcc4),
	.w1(32'hbc1351df),
	.w2(32'hbbaefcca),
	.w3(32'h3c1a1073),
	.w4(32'hbba8edcb),
	.w5(32'h3b8b34ea),
	.w6(32'hbbc6540a),
	.w7(32'hbac1ffe4),
	.w8(32'h3b5a1149),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a2175a),
	.w1(32'hbb4cd5e9),
	.w2(32'h3b83978a),
	.w3(32'h3ab6209f),
	.w4(32'hbbeac6dd),
	.w5(32'h3b3f98be),
	.w6(32'h3b346fc0),
	.w7(32'h3a007175),
	.w8(32'h3b98930b),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a917315),
	.w1(32'hbb09d66d),
	.w2(32'h3afdc8a4),
	.w3(32'hbb351e7c),
	.w4(32'h3bde1826),
	.w5(32'h3ad0f634),
	.w6(32'h3b625eb2),
	.w7(32'h3c1cc8bc),
	.w8(32'h3c37f1d9),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c241f84),
	.w1(32'hbc098d2b),
	.w2(32'hbc33ca6b),
	.w3(32'h3b9a7268),
	.w4(32'hbba60fa3),
	.w5(32'hbcc91229),
	.w6(32'h3c178f74),
	.w7(32'hbbe319a2),
	.w8(32'hbbc75e0f),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a673397),
	.w1(32'hbb99c153),
	.w2(32'hbb6d73b7),
	.w3(32'hbb2e7f01),
	.w4(32'hba1e57c6),
	.w5(32'hbbc7e6ed),
	.w6(32'hbc5a59bb),
	.w7(32'h3b08f9dd),
	.w8(32'h3ab9de63),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb3df0b),
	.w1(32'h3c218965),
	.w2(32'h3be570a0),
	.w3(32'hbad6b293),
	.w4(32'h3b4e7fd5),
	.w5(32'h3cc99725),
	.w6(32'hbb6a7056),
	.w7(32'hbc3e9415),
	.w8(32'hbbed0adb),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2158f2),
	.w1(32'h3a9b7132),
	.w2(32'h3c53c6ea),
	.w3(32'h3b49d780),
	.w4(32'hbbe90442),
	.w5(32'h3c3ca13e),
	.w6(32'hbbe552e8),
	.w7(32'hbc37ed60),
	.w8(32'h39df9506),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baa00b0),
	.w1(32'hbbf01dc0),
	.w2(32'hbc2ed9f5),
	.w3(32'h3b9dbe8f),
	.w4(32'hbc0ecc50),
	.w5(32'hbb88a418),
	.w6(32'h3bc3de50),
	.w7(32'h3c1ee443),
	.w8(32'hbb6a025b),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1245a6),
	.w1(32'hba100aae),
	.w2(32'hbb78a511),
	.w3(32'hbac3c5a0),
	.w4(32'hbbc9938c),
	.w5(32'hba4358c7),
	.w6(32'hbb437131),
	.w7(32'hbb079704),
	.w8(32'h3b033cef),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6c44f3),
	.w1(32'h3ba80952),
	.w2(32'h3c8a3331),
	.w3(32'h3bb0a20a),
	.w4(32'h3a18aa01),
	.w5(32'h3c014b94),
	.w6(32'h3c42bd42),
	.w7(32'h38c97b44),
	.w8(32'hb9cc733d),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbdb07d),
	.w1(32'hbb0f2666),
	.w2(32'h3a9f6cfe),
	.w3(32'h3a40ab72),
	.w4(32'hbc179001),
	.w5(32'hbbb9fb9f),
	.w6(32'h3bafa916),
	.w7(32'hbc1e72d3),
	.w8(32'hbc0dd612),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aef8375),
	.w1(32'h39c4d209),
	.w2(32'hbb99f480),
	.w3(32'h3ba66650),
	.w4(32'h3be7ec62),
	.w5(32'h39b3a684),
	.w6(32'h3bd9facf),
	.w7(32'h3ad574ae),
	.w8(32'hbbcf6da5),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb29a660),
	.w1(32'hbc089c5b),
	.w2(32'hbbf9406c),
	.w3(32'h3a0da35b),
	.w4(32'hbb62a67e),
	.w5(32'hbb9513b9),
	.w6(32'hbbef7a3d),
	.w7(32'h3b84e101),
	.w8(32'hba3e310e),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c10ab58),
	.w1(32'h3c2eb790),
	.w2(32'h3c6c4d31),
	.w3(32'h3b58fa94),
	.w4(32'h3bb15ec0),
	.w5(32'h3c62f379),
	.w6(32'h39564449),
	.w7(32'hba09d10d),
	.w8(32'h3ae56777),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac9d71b),
	.w1(32'h3bd3e5f8),
	.w2(32'h3bd7ddb1),
	.w3(32'hb7a16875),
	.w4(32'h3ac150b5),
	.w5(32'hbb8f7429),
	.w6(32'hba8643ab),
	.w7(32'h3af00b99),
	.w8(32'h3b90209c),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab2ce7d),
	.w1(32'hba92a7f5),
	.w2(32'h3c2fb32c),
	.w3(32'h3b987c87),
	.w4(32'h3a84717c),
	.w5(32'h3b90e91a),
	.w6(32'h3bb7cca5),
	.w7(32'h3c57c534),
	.w8(32'h3c23b96c),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9e3ac2),
	.w1(32'hbb2fae72),
	.w2(32'hbaed52ad),
	.w3(32'hbc1bafd6),
	.w4(32'hbba6d943),
	.w5(32'hbb37c6f5),
	.w6(32'h3ba403b1),
	.w7(32'h3ba72181),
	.w8(32'h3baad8bc),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f0b8d1),
	.w1(32'h3b087aec),
	.w2(32'h3c6f7ede),
	.w3(32'h3bb267f1),
	.w4(32'hbb0098cf),
	.w5(32'hbb21ea55),
	.w6(32'h3b8b870c),
	.w7(32'h3c045239),
	.w8(32'h3ba75b3f),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac82f9c),
	.w1(32'hbb773ac9),
	.w2(32'h3b5eb8cf),
	.w3(32'hbb0724f2),
	.w4(32'h3b44f028),
	.w5(32'hbbcf0974),
	.w6(32'hbb52b8d4),
	.w7(32'hba4f4c81),
	.w8(32'hba826384),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc32dd1b),
	.w1(32'hbbd7481d),
	.w2(32'h3aeecde7),
	.w3(32'hb9ce7e1e),
	.w4(32'hbc036aa5),
	.w5(32'hbc17ae02),
	.w6(32'h3ac3c919),
	.w7(32'hbbe4c91f),
	.w8(32'hbbbd8faf),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb8a727),
	.w1(32'h3beadd7c),
	.w2(32'hbb86ba82),
	.w3(32'hbbd36e6f),
	.w4(32'h3bf54c84),
	.w5(32'hbb934de5),
	.w6(32'h3a86de0c),
	.w7(32'h3b437549),
	.w8(32'hbc4fa326),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfac162),
	.w1(32'hba2a8554),
	.w2(32'h3aedb16e),
	.w3(32'h3bdef62a),
	.w4(32'h3be7be8f),
	.w5(32'h3b274ea3),
	.w6(32'hb925d8de),
	.w7(32'hbba5da82),
	.w8(32'h3a7ed14d),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbda6e36),
	.w1(32'hbba23fb2),
	.w2(32'hbc248dd5),
	.w3(32'hbb8d6166),
	.w4(32'hbb32c2c9),
	.w5(32'hbbb0b1cc),
	.w6(32'hbba26060),
	.w7(32'hbc0662c9),
	.w8(32'hbb56addd),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd0c382),
	.w1(32'hbbf01e1f),
	.w2(32'h3af0170c),
	.w3(32'hbbf04dc3),
	.w4(32'hbba19b63),
	.w5(32'hbb3023aa),
	.w6(32'hbbab891b),
	.w7(32'hb9f47312),
	.w8(32'hb8d6b63b),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba42e69a),
	.w1(32'h3bb15ee8),
	.w2(32'hb9fd2a1c),
	.w3(32'h3ad49999),
	.w4(32'h3b9a56bf),
	.w5(32'h3c81847b),
	.w6(32'h3b87fa19),
	.w7(32'hbc018392),
	.w8(32'h3b319fe7),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc148d8f),
	.w1(32'h3c2221f2),
	.w2(32'h3b093108),
	.w3(32'h3bc22090),
	.w4(32'h3c1ddb85),
	.w5(32'h3893c34e),
	.w6(32'h3bc0e9f1),
	.w7(32'h3b8ccfb3),
	.w8(32'h3b91f5b6),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b633a95),
	.w1(32'h3bd02723),
	.w2(32'hbb7643a9),
	.w3(32'h3c0c8a72),
	.w4(32'h3c440352),
	.w5(32'hbba5bd82),
	.w6(32'h3c179fb6),
	.w7(32'h3ab65e31),
	.w8(32'h3c7ded80),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac9e1bb),
	.w1(32'h3b4ca0a6),
	.w2(32'hb9be5a7f),
	.w3(32'hbc4420ba),
	.w4(32'hbbf19259),
	.w5(32'hbb430578),
	.w6(32'hbc060d8e),
	.w7(32'hbbeb90ee),
	.w8(32'hbbcbf15b),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd46f44),
	.w1(32'h3acfafa1),
	.w2(32'hbc23496d),
	.w3(32'h3c91317f),
	.w4(32'h3c3c233b),
	.w5(32'h3b5e261d),
	.w6(32'h3befcfa0),
	.w7(32'h3b4a87eb),
	.w8(32'h3b912a62),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc50d8bc),
	.w1(32'hbc52e2b8),
	.w2(32'hbc0c5e51),
	.w3(32'hbc18ea42),
	.w4(32'hba9e2f90),
	.w5(32'h3b87f826),
	.w6(32'hbc04480d),
	.w7(32'hbafce0c5),
	.w8(32'hb9152628),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc93163c),
	.w1(32'hbb0b19d6),
	.w2(32'h3aeb4a41),
	.w3(32'hbb64a1f1),
	.w4(32'hbb122a24),
	.w5(32'hbafe47fd),
	.w6(32'hbb196a71),
	.w7(32'hbb0f1e3d),
	.w8(32'hbb831a8d),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb048500),
	.w1(32'hbc2a6177),
	.w2(32'hbc40d4e1),
	.w3(32'hbb4afa98),
	.w4(32'h3b350dc6),
	.w5(32'hbb58f3f6),
	.w6(32'hbc0856cd),
	.w7(32'h3be9b36d),
	.w8(32'hbb802644),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae7aeb7),
	.w1(32'h3b0e4995),
	.w2(32'hbb807178),
	.w3(32'hbb7d7942),
	.w4(32'hbc1d3572),
	.w5(32'hbbb5159a),
	.w6(32'hbba91897),
	.w7(32'hbc0d7544),
	.w8(32'hbb37e44e),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb1929d),
	.w1(32'h3c1f929a),
	.w2(32'h3bfe3f98),
	.w3(32'hbb3c6b98),
	.w4(32'h3b5053e7),
	.w5(32'hbb83f9d1),
	.w6(32'h3be02f07),
	.w7(32'h3bbcd868),
	.w8(32'h3b51c5f9),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c09033e),
	.w1(32'hbc5c6d40),
	.w2(32'hbc4c981b),
	.w3(32'h3ad443f6),
	.w4(32'hbb831873),
	.w5(32'hba6a27a5),
	.w6(32'h3c1b1a5b),
	.w7(32'hbb5fcd35),
	.w8(32'hbc3896bc),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc641c46),
	.w1(32'hbc0f4ca7),
	.w2(32'h3addfd37),
	.w3(32'h3af427d4),
	.w4(32'hb84a26f2),
	.w5(32'hbb81bc5e),
	.w6(32'hbbf57d0f),
	.w7(32'h3be7f1c8),
	.w8(32'h3a9992ef),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c19b491),
	.w1(32'h3aacc0f0),
	.w2(32'h3abe080f),
	.w3(32'h3c0c724a),
	.w4(32'h3bd2fe70),
	.w5(32'hbbe009b6),
	.w6(32'h3c50c2b6),
	.w7(32'h3c28c8e6),
	.w8(32'hbc110973),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc724383),
	.w1(32'hb9ae0a7d),
	.w2(32'h3bb9adf7),
	.w3(32'hbc22811f),
	.w4(32'hbb6a9363),
	.w5(32'hbb5fa524),
	.w6(32'hbc3ec73a),
	.w7(32'hbbb189b2),
	.w8(32'hbc3f015a),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c169ede),
	.w1(32'h3a3f22d9),
	.w2(32'hb91e58ba),
	.w3(32'hba2ff1f1),
	.w4(32'h3b5aa986),
	.w5(32'h3b4aecb7),
	.w6(32'hbae8e91a),
	.w7(32'h3af2cf8d),
	.w8(32'h3b5f201d),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b87fe2b),
	.w1(32'h3af01bf8),
	.w2(32'h3a0b2c1d),
	.w3(32'h3b3d1824),
	.w4(32'h39eeb8ca),
	.w5(32'h35a6936e),
	.w6(32'h3b0ec4e4),
	.w7(32'hba0c434f),
	.w8(32'hba7e7639),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3722c49d),
	.w1(32'h379af845),
	.w2(32'h37d2da1e),
	.w3(32'hb6674807),
	.w4(32'h36a3e46f),
	.w5(32'h378341b4),
	.w6(32'h3717200f),
	.w7(32'h37a7d4cd),
	.w8(32'h380124e4),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b40441c),
	.w1(32'h3b60aabd),
	.w2(32'h3b64ebbf),
	.w3(32'h3aea02bf),
	.w4(32'h3acbc748),
	.w5(32'h3a4faf72),
	.w6(32'h3a8322dc),
	.w7(32'h39f60737),
	.w8(32'h3a440500),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb76d2bb9),
	.w1(32'h3812cc4c),
	.w2(32'h38b55594),
	.w3(32'hb86b1114),
	.w4(32'h36574da8),
	.w5(32'h3820f66d),
	.w6(32'h3824cc25),
	.w7(32'h3891b54a),
	.w8(32'h38e34c10),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af7009b),
	.w1(32'hba85e1f1),
	.w2(32'hb97e485d),
	.w3(32'h3b99c196),
	.w4(32'h3ab157c9),
	.w5(32'h3b25ef68),
	.w6(32'h3b17af79),
	.w7(32'hb9d36c36),
	.w8(32'h3b7225ca),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaae5f54),
	.w1(32'hb8070e2f),
	.w2(32'hba6a4d9e),
	.w3(32'hbb0f60e9),
	.w4(32'hbb05ee5d),
	.w5(32'hbb0f7c03),
	.w6(32'hba10b2aa),
	.w7(32'hba8295bb),
	.w8(32'hba9d1615),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b28effb),
	.w1(32'h3a399e47),
	.w2(32'h389706ae),
	.w3(32'h3ad8120c),
	.w4(32'h3a171094),
	.w5(32'h3843ad86),
	.w6(32'h3b090195),
	.w7(32'h3a0b7877),
	.w8(32'h395ee56d),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396a2b20),
	.w1(32'hb7932e10),
	.w2(32'hba6a43e5),
	.w3(32'hba4f54c8),
	.w4(32'hba85381c),
	.w5(32'hba9b8fa3),
	.w6(32'h380714a9),
	.w7(32'hba0a8623),
	.w8(32'hba907422),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba22352),
	.w1(32'h3b4de75b),
	.w2(32'h3b10d16c),
	.w3(32'h3b852d46),
	.w4(32'h3b2c86e2),
	.w5(32'h3b133bdf),
	.w6(32'h3b63f8d9),
	.w7(32'h3b345c97),
	.w8(32'h3b57d3de),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf90b47),
	.w1(32'h3ba2f1d7),
	.w2(32'h3b8d537f),
	.w3(32'h3bda95ff),
	.w4(32'h3b93e478),
	.w5(32'h3b9ad934),
	.w6(32'h3bb8f59e),
	.w7(32'h3b5d5b36),
	.w8(32'h3b5644de),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca1179b),
	.w1(32'h3a617fd4),
	.w2(32'h3b19c24d),
	.w3(32'h3c92933a),
	.w4(32'h3c1e31be),
	.w5(32'h3c03fb8a),
	.w6(32'h3c59f6a1),
	.w7(32'h3be48449),
	.w8(32'h3bd072b4),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7c221f6),
	.w1(32'hb7d5226d),
	.w2(32'hb7bef7a4),
	.w3(32'h376fff86),
	.w4(32'h384472ed),
	.w5(32'h37f3588e),
	.w6(32'hb7469f55),
	.w7(32'h37a89263),
	.w8(32'hb7c8e489),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94217c1),
	.w1(32'h38964393),
	.w2(32'h399733e7),
	.w3(32'hb8a2a1b9),
	.w4(32'h3900ad97),
	.w5(32'h39a634ee),
	.w6(32'hb962cfa7),
	.w7(32'hb8e2a302),
	.w8(32'h3882cd7d),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa3fc17),
	.w1(32'h3a7b3554),
	.w2(32'h3b4e2a8f),
	.w3(32'hbb877779),
	.w4(32'hbaf03454),
	.w5(32'h3ad1d5f9),
	.w6(32'hba965468),
	.w7(32'hbaacbb46),
	.w8(32'h3abb891d),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd915e3),
	.w1(32'h3c1334fd),
	.w2(32'h3c1822b6),
	.w3(32'h3b35df58),
	.w4(32'h3b5104c9),
	.w5(32'h3b7e5c74),
	.w6(32'h3b598066),
	.w7(32'h3ae3033a),
	.w8(32'h3b8c1162),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be5ddc9),
	.w1(32'h3b62ddbf),
	.w2(32'h3b1234b1),
	.w3(32'h3bc6b4bd),
	.w4(32'h3b3b9bf0),
	.w5(32'h3b02db21),
	.w6(32'h3bc22e31),
	.w7(32'h3b4ada18),
	.w8(32'h3b40dd94),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba25fce3),
	.w1(32'h3ac9ac2e),
	.w2(32'h3acacdbf),
	.w3(32'hba601dfd),
	.w4(32'h3b5837cb),
	.w5(32'h3b8eb754),
	.w6(32'hbba78e6f),
	.w7(32'hbb3e2bb6),
	.w8(32'hbaa419f0),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398579a0),
	.w1(32'h3a210070),
	.w2(32'h3a48f757),
	.w3(32'h38af41ff),
	.w4(32'h39d8773d),
	.w5(32'h39dd71c7),
	.w6(32'h39d991fa),
	.w7(32'h39f1d9c7),
	.w8(32'h39d15dcd),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a26136a),
	.w1(32'h3aaf299c),
	.w2(32'h3ac01e96),
	.w3(32'hb833041f),
	.w4(32'h39b9df31),
	.w5(32'h39c89ed9),
	.w6(32'hb8c7d5e6),
	.w7(32'h38d0b2ea),
	.w8(32'h39559216),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d0f2e),
	.w1(32'hbb895030),
	.w2(32'h3a23d2a4),
	.w3(32'hbb3b4d00),
	.w4(32'hbb99af96),
	.w5(32'hbaced65b),
	.w6(32'hb9885ebd),
	.w7(32'hbb2ebb32),
	.w8(32'hbb73b090),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c541188),
	.w1(32'h3b5aa11e),
	.w2(32'h3c0d3ac4),
	.w3(32'h3c0b3c5d),
	.w4(32'h3b1ebe9c),
	.w5(32'h3b9ea2c1),
	.w6(32'h3b9e8a69),
	.w7(32'hbb656b89),
	.w8(32'h3ae141f1),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b84bb7f),
	.w1(32'hba3e5e35),
	.w2(32'h38d161b8),
	.w3(32'h3b39abd5),
	.w4(32'hb9e17257),
	.w5(32'h3b11093c),
	.w6(32'h3b337b4e),
	.w7(32'h3a18fb52),
	.w8(32'h3a8e30e3),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae514c2),
	.w1(32'hb9bc5cf6),
	.w2(32'hbaafebd5),
	.w3(32'hb98929c3),
	.w4(32'h3a02ffa4),
	.w5(32'hb8b88c9a),
	.w6(32'h39d42307),
	.w7(32'h3ad5355b),
	.w8(32'h3aafa5d4),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc102e7),
	.w1(32'h3bb4df1d),
	.w2(32'h3ba52b0d),
	.w3(32'h3b7e5404),
	.w4(32'h3b6ead69),
	.w5(32'h3b443524),
	.w6(32'h3b039fa7),
	.w7(32'h3b2e5f96),
	.w8(32'h3b1d86e1),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h371484a6),
	.w1(32'h36af08ab),
	.w2(32'h369ec387),
	.w3(32'hb5f6bb65),
	.w4(32'hb6847aee),
	.w5(32'hb62f42c0),
	.w6(32'h37157a47),
	.w7(32'h369c83e2),
	.w8(32'h37047db9),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37919938),
	.w1(32'h371a17a4),
	.w2(32'hb657166c),
	.w3(32'h37024de9),
	.w4(32'hb62b6232),
	.w5(32'hb781339e),
	.w6(32'h369def29),
	.w7(32'hb71227ca),
	.w8(32'hb7386f95),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9d576e),
	.w1(32'h36e0084a),
	.w2(32'hb950765b),
	.w3(32'hba8aaf41),
	.w4(32'h3940c3cc),
	.w5(32'h3a09797d),
	.w6(32'hbaa0952f),
	.w7(32'hb929c0f4),
	.w8(32'h395618fa),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37f063cf),
	.w1(32'h3800ed1a),
	.w2(32'h35bec04c),
	.w3(32'h37ae4dd0),
	.w4(32'h37ee94bf),
	.w5(32'hb6f365d6),
	.w6(32'h38273805),
	.w7(32'h38156e47),
	.w8(32'h379c8eed),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8adc12),
	.w1(32'h3a6eaf34),
	.w2(32'h3afe5a9d),
	.w3(32'hba9a5c95),
	.w4(32'h3a7d084c),
	.w5(32'h3b20e444),
	.w6(32'hbac80841),
	.w7(32'h385b3971),
	.w8(32'h3a339bb1),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb1212f),
	.w1(32'h3c0eb89e),
	.w2(32'h3c193f31),
	.w3(32'h3b12e189),
	.w4(32'h3b259169),
	.w5(32'h3b1344aa),
	.w6(32'h3b65f8e2),
	.w7(32'h3b33386f),
	.w8(32'h3b3786ac),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0bb6e5),
	.w1(32'h3b374568),
	.w2(32'h3b419eb0),
	.w3(32'h3abc5ae9),
	.w4(32'h3b1d674f),
	.w5(32'h3ade029b),
	.w6(32'h3b190054),
	.w7(32'h3abd1310),
	.w8(32'h3aba4c13),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb75a5300),
	.w1(32'hb8118741),
	.w2(32'hb8015689),
	.w3(32'hb78e63a3),
	.w4(32'hb80806dd),
	.w5(32'hb79a9eae),
	.w6(32'hb6ddf76d),
	.w7(32'hb721b7d5),
	.w8(32'h358e7992),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf84318),
	.w1(32'h3b163a68),
	.w2(32'h3b97c607),
	.w3(32'h3bc3aa8f),
	.w4(32'h38bddbd8),
	.w5(32'h3b0a0318),
	.w6(32'h3baa9b21),
	.w7(32'hba646e15),
	.w8(32'hbb5d1786),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b149c2d),
	.w1(32'h3b14cade),
	.w2(32'h3b8ab600),
	.w3(32'h3adeac22),
	.w4(32'h3a83edf9),
	.w5(32'h3b6d6fb0),
	.w6(32'h3b1342cf),
	.w7(32'h3a9d13bf),
	.w8(32'h3b56daf1),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92a7fd4),
	.w1(32'h37a1b64d),
	.w2(32'h39eec45e),
	.w3(32'hb9b96590),
	.w4(32'hb91a03a2),
	.w5(32'h39132f5b),
	.w6(32'hb9c2286e),
	.w7(32'hb9cbf776),
	.w8(32'hb96e5f9f),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b823f4b),
	.w1(32'h3af697f6),
	.w2(32'h3ac7487e),
	.w3(32'h3b5cc8c1),
	.w4(32'h3afd8cfd),
	.w5(32'h3acfd4cc),
	.w6(32'h3b0b0d75),
	.w7(32'h3996f3ac),
	.w8(32'h39628ceb),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3800c7fd),
	.w1(32'h37fd583e),
	.w2(32'h375eaa9e),
	.w3(32'h38402ebe),
	.w4(32'h3809978a),
	.w5(32'h37ca1076),
	.w6(32'h37dd25fa),
	.w7(32'h37774fb1),
	.w8(32'h37db5cfe),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb631ad19),
	.w1(32'h3899e055),
	.w2(32'hb8a72951),
	.w3(32'hb82ab7a9),
	.w4(32'hb87d645f),
	.w5(32'hb983c25d),
	.w6(32'hb8908bc7),
	.w7(32'hb981853b),
	.w8(32'hb9ce11d3),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h383c763e),
	.w1(32'h38489f9d),
	.w2(32'h385d72eb),
	.w3(32'h38068244),
	.w4(32'h37e6f628),
	.w5(32'h37b3296c),
	.w6(32'h36beac63),
	.w7(32'h3601dbb1),
	.w8(32'hb6563f87),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb859cada),
	.w1(32'h361348d1),
	.w2(32'h36882c89),
	.w3(32'hb7c76768),
	.w4(32'h36dc03d4),
	.w5(32'h370e0e44),
	.w6(32'hb6cf8a05),
	.w7(32'h37353fc8),
	.w8(32'h37c042fa),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacb2ab6),
	.w1(32'hbb1674aa),
	.w2(32'hbb54254d),
	.w3(32'hba8ceff5),
	.w4(32'hbb094bd3),
	.w5(32'hbb399695),
	.w6(32'hbb0da950),
	.w7(32'hbadba32d),
	.w8(32'hbb0c40af),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c014296),
	.w1(32'h3bdab7e6),
	.w2(32'h3c37aaa4),
	.w3(32'h3bf9ce3f),
	.w4(32'h3bcbf4d3),
	.w5(32'h3c21a9b4),
	.w6(32'h3ba7b7dd),
	.w7(32'h3b47a266),
	.w8(32'h3bfd1c7b),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bccbc41),
	.w1(32'h3ba9dc1c),
	.w2(32'h3bed970f),
	.w3(32'h3b88cc57),
	.w4(32'h3b0f1659),
	.w5(32'h3b9321be),
	.w6(32'h3b6d72ce),
	.w7(32'h3a33d768),
	.w8(32'h3b333576),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbbc9e5),
	.w1(32'h3b16b8dd),
	.w2(32'h3bbb1b24),
	.w3(32'h3bf10e67),
	.w4(32'h3ba3f477),
	.w5(32'h3bded2e5),
	.w6(32'h3b2f0856),
	.w7(32'h3b306448),
	.w8(32'h3b8784e2),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39432e2e),
	.w1(32'h39852ed9),
	.w2(32'hb83e9e27),
	.w3(32'h3926f01a),
	.w4(32'h3995ddbb),
	.w5(32'h38e7d101),
	.w6(32'h38a60531),
	.w7(32'h39642679),
	.w8(32'h38992e31),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bae180),
	.w1(32'h3a1aa969),
	.w2(32'h3a1431fe),
	.w3(32'h3948a8fb),
	.w4(32'h39937aff),
	.w5(32'h3937d3c4),
	.w6(32'h3820ee28),
	.w7(32'h38fc1a64),
	.w8(32'h3907395a),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36a48526),
	.w1(32'h3519c032),
	.w2(32'hb432afb4),
	.w3(32'hb680087f),
	.w4(32'h37307f54),
	.w5(32'h3696fd86),
	.w6(32'h36dda34f),
	.w7(32'h373834f2),
	.w8(32'h36b550ea),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7dfdae5),
	.w1(32'h36c12b5a),
	.w2(32'hb7b5e3b9),
	.w3(32'h36531959),
	.w4(32'h37325f55),
	.w5(32'hb875693d),
	.w6(32'h37886337),
	.w7(32'hb7e85968),
	.w8(32'hb8b7bc18),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abb5751),
	.w1(32'h3b6b5d7f),
	.w2(32'h3c0b2d27),
	.w3(32'hbaa1fd0e),
	.w4(32'h39703b59),
	.w5(32'h3bb9979b),
	.w6(32'hbb42f777),
	.w7(32'hbb5a17a8),
	.w8(32'h3b96d69b),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37ecb03f),
	.w1(32'h3822c155),
	.w2(32'h380018d3),
	.w3(32'h37cff8a2),
	.w4(32'h3823c9d8),
	.w5(32'h37ce34a8),
	.w6(32'h383abb15),
	.w7(32'h383941b8),
	.w8(32'h37bde298),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6ec6498),
	.w1(32'h3a001c5b),
	.w2(32'hba10a395),
	.w3(32'hba0dc9b1),
	.w4(32'h37c852ab),
	.w5(32'hba11c1ab),
	.w6(32'hba0e6587),
	.w7(32'hba2b3b92),
	.w8(32'hba932dbb),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab33afb),
	.w1(32'h3ab65c1f),
	.w2(32'h3ab10549),
	.w3(32'h3a667c50),
	.w4(32'h3a781830),
	.w5(32'h3a36fb90),
	.w6(32'hb928ac48),
	.w7(32'hb99380c4),
	.w8(32'h38b64f17),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h384be136),
	.w1(32'h3803f18a),
	.w2(32'hb781f9c2),
	.w3(32'h377d9bf0),
	.w4(32'h38067de9),
	.w5(32'hb6059caa),
	.w6(32'h37035977),
	.w7(32'h36dc1bbf),
	.w8(32'hb78f8063),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6a6db9),
	.w1(32'hbae402c1),
	.w2(32'h3ad0fcae),
	.w3(32'h3b0a3c2b),
	.w4(32'hb8fee121),
	.w5(32'h3b03c56f),
	.w6(32'h3b16aab2),
	.w7(32'h39c43f44),
	.w8(32'h3abe782b),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d358aa),
	.w1(32'h3a0f5d7f),
	.w2(32'h3a587158),
	.w3(32'h396bd149),
	.w4(32'h39786166),
	.w5(32'h39dae88b),
	.w6(32'h397f56cd),
	.w7(32'h3998e4f4),
	.w8(32'h39f89fc4),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb7f4b1),
	.w1(32'h3ba8222f),
	.w2(32'h3c3f7ea8),
	.w3(32'h3bbb6f0e),
	.w4(32'h3bc23f79),
	.w5(32'h3c34f019),
	.w6(32'h39a2c492),
	.w7(32'hbaee0e01),
	.w8(32'h3bd4325e),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6ddcabf),
	.w1(32'h38df9ee0),
	.w2(32'h3905574e),
	.w3(32'hb8403669),
	.w4(32'h38c95742),
	.w5(32'h392a175c),
	.w6(32'hb86edf9a),
	.w7(32'h38955736),
	.w8(32'h38ce49d2),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b24681e),
	.w1(32'h3b377491),
	.w2(32'h3b68a52d),
	.w3(32'h3b60ae94),
	.w4(32'h3b56fac9),
	.w5(32'h3bb3f1d2),
	.w6(32'h3b044ad0),
	.w7(32'h39d9cdd7),
	.w8(32'h38fdc998),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule