module layer_10_featuremap_420(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf1d053),
	.w1(32'hbadc4497),
	.w2(32'h3aa8986c),
	.w3(32'hbb4e494d),
	.w4(32'hb90c57aa),
	.w5(32'h39e39f3b),
	.w6(32'hbbe47548),
	.w7(32'h393649e9),
	.w8(32'h38c08b5c),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd9fff9),
	.w1(32'hb75985d0),
	.w2(32'hba8900a1),
	.w3(32'hbb5b714b),
	.w4(32'h39d023ed),
	.w5(32'hbbbf4cbb),
	.w6(32'hbbbc7f1a),
	.w7(32'hbbe6e533),
	.w8(32'hbbe2f83f),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2ab641),
	.w1(32'hbb47eeb5),
	.w2(32'h3b568eb8),
	.w3(32'hba9af7d6),
	.w4(32'hbbbe357c),
	.w5(32'hbbfbed56),
	.w6(32'hbab93425),
	.w7(32'hbaddd461),
	.w8(32'hbb4f6539),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0a0d3c),
	.w1(32'hba1cccc4),
	.w2(32'h3be4a42f),
	.w3(32'hbb96b44a),
	.w4(32'h3b1f180e),
	.w5(32'h3a3e94ab),
	.w6(32'hb9752c40),
	.w7(32'h3b0776e4),
	.w8(32'h3bd29219),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0bf888),
	.w1(32'hbb2fc53b),
	.w2(32'h3ab8b68f),
	.w3(32'h3c1f8b5f),
	.w4(32'h3a973b18),
	.w5(32'hb9806a7c),
	.w6(32'h3ba3000a),
	.w7(32'h39894105),
	.w8(32'hbb1abe91),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9282e3),
	.w1(32'hbb1d5fe6),
	.w2(32'h38d831c1),
	.w3(32'hb98f9caa),
	.w4(32'hbbcc2d9f),
	.w5(32'hbb9ac6bf),
	.w6(32'hb9fe3093),
	.w7(32'hbbaeb7b4),
	.w8(32'hbb1ca9a7),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb93b9ed),
	.w1(32'hbc6857a8),
	.w2(32'hbca3b242),
	.w3(32'hb98664de),
	.w4(32'hbc21b855),
	.w5(32'h3a79d0c3),
	.w6(32'h3ae510dc),
	.w7(32'hb8675682),
	.w8(32'hbc26f47e),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce1c2a6),
	.w1(32'hbcc5191e),
	.w2(32'hbc2395a7),
	.w3(32'hbc974c7f),
	.w4(32'hbc7807bb),
	.w5(32'hbbe3156f),
	.w6(32'hbcab8566),
	.w7(32'hbc53ee43),
	.w8(32'hbb885ac5),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ec56e0),
	.w1(32'hbb4316cd),
	.w2(32'hbac87843),
	.w3(32'hb9608877),
	.w4(32'hbb972eac),
	.w5(32'hbbce8c76),
	.w6(32'h3aa4ba78),
	.w7(32'h39276174),
	.w8(32'hbb1ac07a),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc63d8d6),
	.w1(32'hbc1da998),
	.w2(32'hbcaf01ed),
	.w3(32'h3ac1aed4),
	.w4(32'h3aca6c61),
	.w5(32'hbc004e24),
	.w6(32'hbbd228a2),
	.w7(32'hbb587dab),
	.w8(32'hbc01ed02),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb09dffa),
	.w1(32'h3b606fb7),
	.w2(32'h3a7a0d47),
	.w3(32'h3bc2f65a),
	.w4(32'h3b1aa207),
	.w5(32'h3951e1fa),
	.w6(32'h3a850257),
	.w7(32'h3a598ed5),
	.w8(32'h3a2e7431),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb983e8d8),
	.w1(32'hbbb12f27),
	.w2(32'hbc53274d),
	.w3(32'h3bf7eecb),
	.w4(32'hbbadffaf),
	.w5(32'hbbf20274),
	.w6(32'hbad0aea6),
	.w7(32'h39768723),
	.w8(32'hbbf2d5b8),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb88fc65),
	.w1(32'hbb18a332),
	.w2(32'hbc37895c),
	.w3(32'h3c095951),
	.w4(32'h3c3fe42f),
	.w5(32'hbb908dd8),
	.w6(32'h3bd2a17a),
	.w7(32'hba7669b7),
	.w8(32'hbbd296ca),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7df286),
	.w1(32'hbc1bc330),
	.w2(32'hbc534717),
	.w3(32'h3b7bb175),
	.w4(32'hbb877cf6),
	.w5(32'hbc4a53dc),
	.w6(32'h3ae6bd4f),
	.w7(32'hbac11223),
	.w8(32'hbc09486f),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba1f2e0),
	.w1(32'hbb219d7b),
	.w2(32'hba0057e0),
	.w3(32'hbb38c40e),
	.w4(32'h3b9d8928),
	.w5(32'hbb7a6832),
	.w6(32'hbb05eb9b),
	.w7(32'h3a4ee761),
	.w8(32'hbbbac426),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3d1af0),
	.w1(32'hbc5570a9),
	.w2(32'hbc5b423b),
	.w3(32'hbc671cdd),
	.w4(32'h3a1fe429),
	.w5(32'h3b1a75db),
	.w6(32'hbc89e465),
	.w7(32'hbbeed796),
	.w8(32'hbc77fbc9),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9f9c64),
	.w1(32'h3a8f0c22),
	.w2(32'h3b192087),
	.w3(32'hb926baec),
	.w4(32'h3b358ee3),
	.w5(32'h3ae40996),
	.w6(32'h3acd7cab),
	.w7(32'h3b596600),
	.w8(32'h3bd33302),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc854c78),
	.w1(32'hbc4c04ea),
	.w2(32'hbcaa9fd3),
	.w3(32'hbc003467),
	.w4(32'h392b7776),
	.w5(32'hbc397451),
	.w6(32'hbc1b8eeb),
	.w7(32'hbb8efc95),
	.w8(32'hbc962968),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0eb0a3),
	.w1(32'hba9a3267),
	.w2(32'hbbc898b3),
	.w3(32'hba319e8f),
	.w4(32'h3a92a2c7),
	.w5(32'h3b197e94),
	.w6(32'hbb3e15ce),
	.w7(32'h3ab0c7ba),
	.w8(32'hbbd42235),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1b9671),
	.w1(32'h3b0973a6),
	.w2(32'hbb8269e3),
	.w3(32'h3b645ada),
	.w4(32'hba79660c),
	.w5(32'hbba33db7),
	.w6(32'h3b51ea53),
	.w7(32'hba5aadcc),
	.w8(32'hba40a5f7),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b02fad5),
	.w1(32'hb96ad33c),
	.w2(32'hbb7020fe),
	.w3(32'h3a8a600e),
	.w4(32'hbb64ad05),
	.w5(32'hbbd96117),
	.w6(32'hbaf9924d),
	.w7(32'hbb349441),
	.w8(32'hbbbe61a1),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaad6519),
	.w1(32'h3b0c6093),
	.w2(32'h37e42af8),
	.w3(32'hbb8bfe66),
	.w4(32'h3a5adcda),
	.w5(32'hbb158320),
	.w6(32'h3a00c521),
	.w7(32'h3b73d68a),
	.w8(32'hba36b889),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca8a85f),
	.w1(32'hbcb8bdc1),
	.w2(32'hbd084513),
	.w3(32'hbbf0099b),
	.w4(32'hba84895f),
	.w5(32'hbb3b784f),
	.w6(32'hbd0cfb06),
	.w7(32'hbc623f04),
	.w8(32'hbd090aad),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb60366c),
	.w1(32'hbb5dac96),
	.w2(32'hbc7cd927),
	.w3(32'h3b907108),
	.w4(32'h3b8a657e),
	.w5(32'hbbeee875),
	.w6(32'hbbf037f3),
	.w7(32'hbbaed5b2),
	.w8(32'hbc9ae497),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb700ea7),
	.w1(32'h3be03d77),
	.w2(32'hbae98c8e),
	.w3(32'hbc098597),
	.w4(32'h3c029d1c),
	.w5(32'hbbc32636),
	.w6(32'hbc5472f5),
	.w7(32'hbbb01918),
	.w8(32'hbc59c02c),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5799a7),
	.w1(32'h3afd7053),
	.w2(32'h3b11da9e),
	.w3(32'hba0c5a63),
	.w4(32'h398c6390),
	.w5(32'h39f00538),
	.w6(32'hbb1f2880),
	.w7(32'h3b883786),
	.w8(32'h3b70fef8),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abd07ee),
	.w1(32'h3a94f485),
	.w2(32'h3a1949af),
	.w3(32'h39f9a823),
	.w4(32'h3b1997de),
	.w5(32'h3b355166),
	.w6(32'h3bdbbefd),
	.w7(32'h3b44c8fd),
	.w8(32'hbb3a104e),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ccaea2f),
	.w1(32'hbc6610b3),
	.w2(32'hbc812c73),
	.w3(32'h3c5116ec),
	.w4(32'hbc49f876),
	.w5(32'hb9723721),
	.w6(32'h3cd7639b),
	.w7(32'hbb14187d),
	.w8(32'hbbe3cfb2),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6c842d),
	.w1(32'h39c28551),
	.w2(32'h3b14ffd6),
	.w3(32'hba593484),
	.w4(32'hbab7b704),
	.w5(32'h3b59146a),
	.w6(32'hbb223f2e),
	.w7(32'h3aed4ffd),
	.w8(32'h3b021ff5),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce1cfeb),
	.w1(32'h3bd8db88),
	.w2(32'hbb22039e),
	.w3(32'h3c200630),
	.w4(32'hbb44684e),
	.w5(32'hbc6ae8d9),
	.w6(32'h3c009674),
	.w7(32'hbc58ad90),
	.w8(32'hbcb32905),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb62abfd),
	.w1(32'h3bddb84a),
	.w2(32'h3ac40f39),
	.w3(32'hbb996c4a),
	.w4(32'h3b1de4dc),
	.w5(32'h3aedcb63),
	.w6(32'hbb891028),
	.w7(32'h389ff6a5),
	.w8(32'h3b5d339e),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37c12e80),
	.w1(32'h3aed8519),
	.w2(32'h38fe4b3f),
	.w3(32'hbb2e409f),
	.w4(32'h39d44d04),
	.w5(32'hbb9e70c5),
	.w6(32'h3b1b95b9),
	.w7(32'h3a7428b1),
	.w8(32'hba4b93de),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb95fd51),
	.w1(32'hbadffff3),
	.w2(32'hbc09bbe9),
	.w3(32'hbad494ba),
	.w4(32'h3b585059),
	.w5(32'hbbcee922),
	.w6(32'hbb5fdfb5),
	.w7(32'hba42aa8d),
	.w8(32'hbb6788da),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb45489a),
	.w1(32'hbb139065),
	.w2(32'hbbec1d76),
	.w3(32'hbbe61d01),
	.w4(32'hbb5488d5),
	.w5(32'h3b7a08c5),
	.w6(32'hbabf1fdd),
	.w7(32'hbba50c67),
	.w8(32'hbb9f2713),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9259e7),
	.w1(32'h3aaaaf96),
	.w2(32'hbbd18f72),
	.w3(32'hbb0ec4a8),
	.w4(32'hb9a168b3),
	.w5(32'hbb200a39),
	.w6(32'hba83e4dc),
	.w7(32'hb9d2230c),
	.w8(32'hba02d78d),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8533bc),
	.w1(32'hbc2c2d1c),
	.w2(32'hbc21bd07),
	.w3(32'h3b05450e),
	.w4(32'hbbe214a6),
	.w5(32'hbc2f5342),
	.w6(32'h3b75582f),
	.w7(32'hb9f33c53),
	.w8(32'hbadb620d),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcdf31de),
	.w1(32'hbc3c9f21),
	.w2(32'hbc96e121),
	.w3(32'h3af14b7f),
	.w4(32'h3c0652c8),
	.w5(32'h3be10121),
	.w6(32'hbc32eb8b),
	.w7(32'h3c04ec3b),
	.w8(32'h3b3e7669),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c68f524),
	.w1(32'h3c587275),
	.w2(32'hbb0dfdaa),
	.w3(32'h3c2749a5),
	.w4(32'h3c4d96cb),
	.w5(32'hbbe72d98),
	.w6(32'hbafc20c1),
	.w7(32'hbc07d53a),
	.w8(32'hbc544d43),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cfb5b7c),
	.w1(32'hbb2ae631),
	.w2(32'hbcac8c7e),
	.w3(32'h3ca1cd5f),
	.w4(32'hbc02d2fc),
	.w5(32'hbcd01dfd),
	.w6(32'h3c9fc39a),
	.w7(32'hbc2eef3f),
	.w8(32'hbcf6a7ba),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac9c1c7),
	.w1(32'h3b1c15c7),
	.w2(32'h3aae68b2),
	.w3(32'h3ab5d2a8),
	.w4(32'h393f1d88),
	.w5(32'hbac030f1),
	.w6(32'hbad0dac9),
	.w7(32'hbadbc720),
	.w8(32'hba0b40b8),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2067a4),
	.w1(32'hbb807431),
	.w2(32'h3adfa015),
	.w3(32'h3a9f2376),
	.w4(32'h3c077b39),
	.w5(32'hb95d10df),
	.w6(32'h3b255d1f),
	.w7(32'h3a7b007b),
	.w8(32'hbb562dc8),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4695c1),
	.w1(32'hbb54914a),
	.w2(32'h3a8675df),
	.w3(32'h3a9d1a77),
	.w4(32'h39c31796),
	.w5(32'h3c4568af),
	.w6(32'hb992d761),
	.w7(32'h3836ce19),
	.w8(32'h3b62f8d3),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399a40d3),
	.w1(32'h3b1ccd7e),
	.w2(32'h3bc7284c),
	.w3(32'hbbc1d0b0),
	.w4(32'h3be11bb6),
	.w5(32'hbac78f4c),
	.w6(32'hbb47a5f7),
	.w7(32'h3b560ff2),
	.w8(32'h3b83d6e7),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc806b1d),
	.w1(32'hbc4809f2),
	.w2(32'hbcbcf0e4),
	.w3(32'hbb5d33e4),
	.w4(32'h3a9eef44),
	.w5(32'hbbab69f0),
	.w6(32'hbbcecc2d),
	.w7(32'hb9a953c7),
	.w8(32'hbc6835c9),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ee8da),
	.w1(32'h3a6d36d5),
	.w2(32'hbbb1537e),
	.w3(32'hbac8fe4e),
	.w4(32'h3bad3743),
	.w5(32'h3bb34ad7),
	.w6(32'hbbf0441e),
	.w7(32'hbb839d8b),
	.w8(32'hbc366c49),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbba1142),
	.w1(32'hbb35694a),
	.w2(32'hbc36a503),
	.w3(32'h3bb1fb19),
	.w4(32'h3c4b152f),
	.w5(32'h3b42f79d),
	.w6(32'hbc484966),
	.w7(32'hbb86c5ed),
	.w8(32'hbc6eba4f),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfed5c1),
	.w1(32'hbb48be5d),
	.w2(32'hbbab60db),
	.w3(32'hbb3fc7a8),
	.w4(32'h3bffc3f3),
	.w5(32'hbbd84f4a),
	.w6(32'hbc19c7bd),
	.w7(32'hbba926d7),
	.w8(32'hbc80fcfe),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1a9071),
	.w1(32'hbc27bc38),
	.w2(32'hbcc49da3),
	.w3(32'h3c0a655f),
	.w4(32'h3b35b50e),
	.w5(32'hbc18f603),
	.w6(32'hbc023893),
	.w7(32'hbb7382de),
	.w8(32'hbca66066),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac53287),
	.w1(32'h3ae9a8dd),
	.w2(32'hb9d216c6),
	.w3(32'hbaed0afa),
	.w4(32'hbb307411),
	.w5(32'hbb422789),
	.w6(32'hbb838155),
	.w7(32'h3b329ef2),
	.w8(32'hba735394),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa659e5),
	.w1(32'hbb75a36d),
	.w2(32'hba256192),
	.w3(32'hbb09698a),
	.w4(32'hbb59be5c),
	.w5(32'h3a452729),
	.w6(32'h3b58a76b),
	.w7(32'hba674541),
	.w8(32'hbaae3ad8),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dc3aa8),
	.w1(32'h3a0c8fd2),
	.w2(32'h3b46ede7),
	.w3(32'hbb81daf2),
	.w4(32'hbb56632f),
	.w5(32'h3b68826b),
	.w6(32'h3baaec13),
	.w7(32'h39da6f2b),
	.w8(32'h3a440260),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbed4037),
	.w1(32'hbbb9c101),
	.w2(32'hbc5ea287),
	.w3(32'hbbb576ba),
	.w4(32'hba9c2897),
	.w5(32'hbc15feb8),
	.w6(32'hbb99a78d),
	.w7(32'hbabcfceb),
	.w8(32'hbc2581c0),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb22da32),
	.w1(32'hb9f5cb80),
	.w2(32'hbb49dea4),
	.w3(32'h39dba953),
	.w4(32'hba947403),
	.w5(32'h3b942d53),
	.w6(32'hbaa40dca),
	.w7(32'hbb09e274),
	.w8(32'hbb3f9bad),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc835334),
	.w1(32'hbbd21ed7),
	.w2(32'hbcb0aafd),
	.w3(32'hbb28f07e),
	.w4(32'hb9debf31),
	.w5(32'hbc45884a),
	.w6(32'hbbbd070c),
	.w7(32'hbb61ecb3),
	.w8(32'hbc8f3d6c),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb268dd9),
	.w1(32'hbb89fcd9),
	.w2(32'hbc15abff),
	.w3(32'hbb8ffb65),
	.w4(32'hbba87393),
	.w5(32'hbc392401),
	.w6(32'h3a971b67),
	.w7(32'hbc03725c),
	.w8(32'hbb2bec0a),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f09963),
	.w1(32'hb9513af9),
	.w2(32'hbb12f326),
	.w3(32'hbace2833),
	.w4(32'h3a7af878),
	.w5(32'hbc3396f1),
	.w6(32'h39030c45),
	.w7(32'hbb07aa02),
	.w8(32'h3b871960),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb842406),
	.w1(32'h3a991c8f),
	.w2(32'h3b46e1e4),
	.w3(32'h39e08b0d),
	.w4(32'h3bb70601),
	.w5(32'h3bc379ae),
	.w6(32'h3b82c318),
	.w7(32'h3aeef86a),
	.w8(32'h3b0f6113),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb89e97),
	.w1(32'hbac7e26e),
	.w2(32'hbac24a33),
	.w3(32'h3b7cbeac),
	.w4(32'hbb07567e),
	.w5(32'hbb3bd898),
	.w6(32'h3acabdca),
	.w7(32'hb8f7d393),
	.w8(32'hbbadcf90),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9b3486),
	.w1(32'h3a9637c0),
	.w2(32'h3ab3ad5a),
	.w3(32'h3a9ea8cf),
	.w4(32'hb91a09e0),
	.w5(32'h3b94f764),
	.w6(32'h3b7a2a6c),
	.w7(32'h3bbc0c90),
	.w8(32'h3b296e78),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac38396),
	.w1(32'h3ad0ec91),
	.w2(32'h37a6cf8b),
	.w3(32'hbb729f93),
	.w4(32'hb9c331a0),
	.w5(32'hbbcc5f2e),
	.w6(32'hbb863f95),
	.w7(32'h3abd0633),
	.w8(32'hbb29631c),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc279881),
	.w1(32'hbb21ceab),
	.w2(32'hbc140872),
	.w3(32'h3a04f521),
	.w4(32'hbb3b9796),
	.w5(32'hbbacf3a7),
	.w6(32'hbb5af61a),
	.w7(32'hbb52fc84),
	.w8(32'hbbeb4e89),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1a95e8),
	.w1(32'hbc16b1b8),
	.w2(32'hbc05500f),
	.w3(32'hbc129a55),
	.w4(32'hbbd1258c),
	.w5(32'hbb9124fe),
	.w6(32'hba9e25c4),
	.w7(32'h3b9e1114),
	.w8(32'hbb9e9a0d),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9a2a40),
	.w1(32'hbb82bb16),
	.w2(32'h3ac87712),
	.w3(32'hbb0f3dd5),
	.w4(32'h3b65a4f7),
	.w5(32'hbb1c7369),
	.w6(32'h39d25fce),
	.w7(32'hbaa1623c),
	.w8(32'h3adb5cc4),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0395f6),
	.w1(32'hbab622f1),
	.w2(32'h3b3f313c),
	.w3(32'h3baed329),
	.w4(32'hb79eeecf),
	.w5(32'h3bb0c642),
	.w6(32'h3adfc5af),
	.w7(32'h3a4a0ece),
	.w8(32'hba6765fd),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9da905a),
	.w1(32'h3b9781f0),
	.w2(32'h3b392040),
	.w3(32'h3b30c137),
	.w4(32'h3b827ce3),
	.w5(32'hbb850b57),
	.w6(32'h3af0a9c2),
	.w7(32'h3afb5d1a),
	.w8(32'hb96cd5de),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3408f2),
	.w1(32'hbadf6b3b),
	.w2(32'hba85f3c5),
	.w3(32'h3b98f2dd),
	.w4(32'hbb00557d),
	.w5(32'h3c005c6c),
	.w6(32'h3befc8ef),
	.w7(32'h39ed68fd),
	.w8(32'h3b1b76a4),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca9216e),
	.w1(32'hbc77bdfb),
	.w2(32'hbc9cc73e),
	.w3(32'h3a89c893),
	.w4(32'hbb536179),
	.w5(32'hbb70203c),
	.w6(32'hbbe96740),
	.w7(32'hbb4b925c),
	.w8(32'hbc61290f),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcc1b4d),
	.w1(32'hbc0f31d0),
	.w2(32'hbca372de),
	.w3(32'h3c09e056),
	.w4(32'h3b28ec6c),
	.w5(32'hbba74bd5),
	.w6(32'hbcd38f04),
	.w7(32'hbc874d01),
	.w8(32'hbc927311),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7eb85c),
	.w1(32'hbc4754f1),
	.w2(32'hbcadd3a4),
	.w3(32'hbc4a6260),
	.w4(32'hbae71e57),
	.w5(32'hbc8903fd),
	.w6(32'hbc88d60c),
	.w7(32'hbbcba04b),
	.w8(32'hbca14ab5),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdd8077),
	.w1(32'h3b41f5be),
	.w2(32'hbc6fe151),
	.w3(32'h3b2af9f8),
	.w4(32'h3b98c2b3),
	.w5(32'hbbe2a719),
	.w6(32'hbc2f5df9),
	.w7(32'hbc8570e0),
	.w8(32'hbd045e2d),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc049fca),
	.w1(32'h3b07cce7),
	.w2(32'h3b97bb62),
	.w3(32'hbc26f3cc),
	.w4(32'h3b117371),
	.w5(32'h3bd07775),
	.w6(32'hbc22c6ef),
	.w7(32'h3b873b98),
	.w8(32'h3ac37454),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b80d86e),
	.w1(32'hbabbf660),
	.w2(32'h38d60687),
	.w3(32'hb7b41d24),
	.w4(32'h398030bb),
	.w5(32'h3b1caad6),
	.w6(32'hbb8e9509),
	.w7(32'h3b4e2e4a),
	.w8(32'h3bcf7250),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b60ec52),
	.w1(32'hb8c74f56),
	.w2(32'h3a6883fe),
	.w3(32'h3c37f87f),
	.w4(32'h3b54d2c1),
	.w5(32'h3be999bf),
	.w6(32'h3b2fd87e),
	.w7(32'h3bbaeaa8),
	.w8(32'h3b1cbcc6),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ac168),
	.w1(32'hbb3c2c17),
	.w2(32'hbb77c130),
	.w3(32'hbbab2b77),
	.w4(32'h3afe9d83),
	.w5(32'hbbbfa451),
	.w6(32'hbbbecb20),
	.w7(32'hb9d43e86),
	.w8(32'hbbdf3f29),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb097554),
	.w1(32'h3bc2818f),
	.w2(32'h3b6fdb9d),
	.w3(32'hbba09930),
	.w4(32'h3a98d8f9),
	.w5(32'hbb556b6b),
	.w6(32'hbb81ede2),
	.w7(32'h3bbc9bfe),
	.w8(32'h3b955f8b),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc744a4e),
	.w1(32'hbbb5d1bb),
	.w2(32'hbbd05c8c),
	.w3(32'hbbb645c2),
	.w4(32'hbbdbbd07),
	.w5(32'hbb3165ae),
	.w6(32'h3b926e34),
	.w7(32'hba9c22a6),
	.w8(32'hbb1a1ca1),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc38bd6e),
	.w1(32'hbbd2a607),
	.w2(32'hbc814ef1),
	.w3(32'h3b0d218f),
	.w4(32'h3b81646f),
	.w5(32'hbbade563),
	.w6(32'hbc1346f6),
	.w7(32'h38faf0a2),
	.w8(32'hbc39a10c),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc25a232),
	.w1(32'hbab591f9),
	.w2(32'hbbb62679),
	.w3(32'h3a01fc6f),
	.w4(32'h3bb3e998),
	.w5(32'h3bfe3b5a),
	.w6(32'hbc019dc4),
	.w7(32'hbbd27293),
	.w8(32'hbb8de1eb),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9184e1),
	.w1(32'hbb84fc2c),
	.w2(32'hbb2012e3),
	.w3(32'hba8e6d46),
	.w4(32'hbb2e58f7),
	.w5(32'h3ba3c6c8),
	.w6(32'hbbbf531f),
	.w7(32'hbba372db),
	.w8(32'hbb19cfbf),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc11ef24),
	.w1(32'hbbd1b35c),
	.w2(32'hbc3a4de8),
	.w3(32'h3be02ab4),
	.w4(32'hbb391f1f),
	.w5(32'hbbcab1d1),
	.w6(32'hb89ba294),
	.w7(32'h3a15da1d),
	.w8(32'hbc331eef),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2401b5),
	.w1(32'h3b9e8bd1),
	.w2(32'hbacabde3),
	.w3(32'hbc090ca0),
	.w4(32'h3bf8be1b),
	.w5(32'h3a939013),
	.w6(32'hbc036257),
	.w7(32'h3b60b190),
	.w8(32'hbb65c637),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc14ed21),
	.w1(32'hba1be215),
	.w2(32'hbc142588),
	.w3(32'hbbcec33a),
	.w4(32'h39e8d276),
	.w5(32'hbb6cc30e),
	.w6(32'hbc343cc2),
	.w7(32'hb920a005),
	.w8(32'hbbe3a6d3),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac9a0e1),
	.w1(32'h3ae73386),
	.w2(32'h39803064),
	.w3(32'h3b2d5dec),
	.w4(32'h3b366b15),
	.w5(32'h3a8f766f),
	.w6(32'h3b32b430),
	.w7(32'h3a8259b3),
	.w8(32'h3b0386e9),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b125fe3),
	.w1(32'hbc134c21),
	.w2(32'hbbce7765),
	.w3(32'h38cf42ed),
	.w4(32'hbb9f42e5),
	.w5(32'hbbd595ef),
	.w6(32'hbb8ed18c),
	.w7(32'hbbc5439d),
	.w8(32'hbbefda0d),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc329b67),
	.w1(32'h3bce04f3),
	.w2(32'h3a9355c1),
	.w3(32'hbc530909),
	.w4(32'h3b370f2c),
	.w5(32'h3bab5155),
	.w6(32'hbb7ebb07),
	.w7(32'h3bbe9637),
	.w8(32'h3ba7004c),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb00f9bf),
	.w1(32'hbb19ff8a),
	.w2(32'h3af8bdaf),
	.w3(32'hbaeaf4f7),
	.w4(32'hbbd21501),
	.w5(32'hbb95bc84),
	.w6(32'h3a70dba1),
	.w7(32'hbb93f5a2),
	.w8(32'hb9c4466f),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abd4ab0),
	.w1(32'h3b2a15f7),
	.w2(32'h3ae684b4),
	.w3(32'h3b93d968),
	.w4(32'h3b87c80b),
	.w5(32'h3bf61142),
	.w6(32'h3b258b43),
	.w7(32'hbb663d49),
	.w8(32'hbbea40a6),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1940e0),
	.w1(32'hbb3eb938),
	.w2(32'hb997d1af),
	.w3(32'h3bcc45c3),
	.w4(32'hbb0b792d),
	.w5(32'hbacc4335),
	.w6(32'h3b913cdb),
	.w7(32'h3aff6517),
	.w8(32'h3bdb8625),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb186dfb),
	.w1(32'h3aa16bbf),
	.w2(32'h3b612aa1),
	.w3(32'h3b6cd0b0),
	.w4(32'h3bd71480),
	.w5(32'h3b8564cf),
	.w6(32'h3ab311cb),
	.w7(32'hbbe49ded),
	.w8(32'hbc210f68),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9a9451),
	.w1(32'hbc169083),
	.w2(32'hbc75732d),
	.w3(32'hbc18d90c),
	.w4(32'hbb5ea41c),
	.w5(32'hbbcb8627),
	.w6(32'hbcc3cc57),
	.w7(32'hbc605dbe),
	.w8(32'hbcbc7d1f),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c90ab58),
	.w1(32'h3b828f86),
	.w2(32'hb756e178),
	.w3(32'h3c4a7ca7),
	.w4(32'hbb493875),
	.w5(32'hbb3e8efb),
	.w6(32'h3c635d86),
	.w7(32'hbbf461d2),
	.w8(32'hbbf5bdc3),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8c9f5a),
	.w1(32'hbc3d8516),
	.w2(32'hbc65bd07),
	.w3(32'hb7c9f83c),
	.w4(32'hbb3df280),
	.w5(32'hbb80f7b2),
	.w6(32'hbc7c65da),
	.w7(32'hbaf3671d),
	.w8(32'hbc38dbe4),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb50e41),
	.w1(32'h3b59c694),
	.w2(32'hbb28ff3b),
	.w3(32'hbb795c6a),
	.w4(32'hbb7c5b2e),
	.w5(32'hbc03f579),
	.w6(32'hba500221),
	.w7(32'hbc253bcc),
	.w8(32'hbc0fa905),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc93dc66),
	.w1(32'hbbc717f6),
	.w2(32'hbbe23ae0),
	.w3(32'hbbc469a4),
	.w4(32'h3ba9c5d7),
	.w5(32'h3b977a30),
	.w6(32'hbc991f73),
	.w7(32'hbc301509),
	.w8(32'hbc3a0af6),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba6c4c6),
	.w1(32'hbbc0e6e6),
	.w2(32'hbab16cea),
	.w3(32'hbb05089a),
	.w4(32'hbb4ccb2d),
	.w5(32'hbc024eeb),
	.w6(32'hbba80bdc),
	.w7(32'hbb557989),
	.w8(32'hbc1cb7e6),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9a637f),
	.w1(32'hbc0c5373),
	.w2(32'hbb9a3bf5),
	.w3(32'hbae53ded),
	.w4(32'hba5e4ee7),
	.w5(32'hbb0b69c6),
	.w6(32'h3bdee29b),
	.w7(32'hbc123444),
	.w8(32'hbbd3f07e),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbce92c1),
	.w1(32'hbb63f834),
	.w2(32'hbb46535e),
	.w3(32'hbbcc4311),
	.w4(32'hbb82cea8),
	.w5(32'hba250f4f),
	.w6(32'h3b09e7d1),
	.w7(32'h3a172c9c),
	.w8(32'h3a97f780),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb964476),
	.w1(32'hbbc40c24),
	.w2(32'hbc843d6e),
	.w3(32'h3ae2106b),
	.w4(32'h3b4cc3c4),
	.w5(32'hbbe008d7),
	.w6(32'hbbb99289),
	.w7(32'hbb125ede),
	.w8(32'hbcafb0a6),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2a1c26),
	.w1(32'hbc254efb),
	.w2(32'hbc9d71bf),
	.w3(32'h3982a254),
	.w4(32'hbc094be1),
	.w5(32'hbc6fd974),
	.w6(32'hbb823fcb),
	.w7(32'hbc18b168),
	.w8(32'hbca593ea),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce61a5d),
	.w1(32'hbc94fb04),
	.w2(32'hbce47cb2),
	.w3(32'hbc80b9b0),
	.w4(32'hbb5f21fe),
	.w5(32'hba90d59b),
	.w6(32'hbd24e3ef),
	.w7(32'hbaca4248),
	.w8(32'hbc1a0e66),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba10bef8),
	.w1(32'h3bd7cb07),
	.w2(32'h3bceba4d),
	.w3(32'hbb64fc74),
	.w4(32'h3c0a7d15),
	.w5(32'h3c0e66f3),
	.w6(32'hbc4ac66c),
	.w7(32'h3aba6f77),
	.w8(32'hbb0025a5),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1668d7),
	.w1(32'hbb9ae17c),
	.w2(32'hbc1c45ed),
	.w3(32'h3b82ec65),
	.w4(32'hbb15c89a),
	.w5(32'h38fe4e33),
	.w6(32'hbc01ca65),
	.w7(32'hbc6ab8c1),
	.w8(32'hbc47e1bb),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc900171),
	.w1(32'hbc9306bd),
	.w2(32'hbcb55137),
	.w3(32'h3b534183),
	.w4(32'hbb2b51c7),
	.w5(32'hbb3a891c),
	.w6(32'hbbf7eb60),
	.w7(32'h3bc3904b),
	.w8(32'hbbe5267c),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb728510),
	.w1(32'h3bc9bb1e),
	.w2(32'h3c07e1e5),
	.w3(32'hbb1c4846),
	.w4(32'h3b43268a),
	.w5(32'h3c594624),
	.w6(32'h3b2201f5),
	.w7(32'h3ba1e616),
	.w8(32'h3c215029),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcfdc93b),
	.w1(32'hbc85637b),
	.w2(32'hbcaaaf25),
	.w3(32'hbbd0b760),
	.w4(32'hbb93975d),
	.w5(32'hbc5498b5),
	.w6(32'hbc6f8715),
	.w7(32'hbbc4ca81),
	.w8(32'hbc38d5ef),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb09f183),
	.w1(32'hbbc06e5a),
	.w2(32'hbc8c88f6),
	.w3(32'h3ba58a14),
	.w4(32'hbc0abfa6),
	.w5(32'hbca2f7e1),
	.w6(32'hbac45228),
	.w7(32'hbba4527d),
	.w8(32'hbc32c82a),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4ba6d0),
	.w1(32'h3bd6932e),
	.w2(32'h3b5bf4a4),
	.w3(32'hbbbf9c5d),
	.w4(32'h3ba1d59e),
	.w5(32'h3c00ab84),
	.w6(32'hbb8a9f31),
	.w7(32'h3b364b5a),
	.w8(32'h3bbbd13c),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5f85f3a),
	.w1(32'hbb9c2a7e),
	.w2(32'hbbd675b3),
	.w3(32'h3aed8cd6),
	.w4(32'hbb2f1d04),
	.w5(32'h3b2de92b),
	.w6(32'h3aa4ec58),
	.w7(32'hbbc17be8),
	.w8(32'hbb952c6a),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb944b02),
	.w1(32'h3aa84f70),
	.w2(32'hbc1e09f3),
	.w3(32'h3a690dfb),
	.w4(32'h3bd53189),
	.w5(32'hbbe16c3b),
	.w6(32'hbb79e418),
	.w7(32'hbb035c81),
	.w8(32'hbc4c60fa),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdf18b0),
	.w1(32'hbb5aa746),
	.w2(32'hbc119bf8),
	.w3(32'h3bb2bd44),
	.w4(32'hba6786e7),
	.w5(32'hbbd93425),
	.w6(32'hbae6f429),
	.w7(32'hbb9681d0),
	.w8(32'hbc2974f3),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6b846f),
	.w1(32'hb8d4b544),
	.w2(32'hbbb0a99e),
	.w3(32'h3b8dc3d4),
	.w4(32'h3ae51643),
	.w5(32'h3abd50df),
	.w6(32'h3b60ea66),
	.w7(32'h3b0d528e),
	.w8(32'hbaa7d65b),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb46cf5e),
	.w1(32'hbb82b98b),
	.w2(32'hbbb8db74),
	.w3(32'h3b551c70),
	.w4(32'hbadf50bf),
	.w5(32'hbb872ffa),
	.w6(32'h3bbc50a3),
	.w7(32'hbbf1c1bc),
	.w8(32'hbc60e0e4),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb45e25),
	.w1(32'hb98b3717),
	.w2(32'h39f9217d),
	.w3(32'h3b3ac23b),
	.w4(32'h3ba159ac),
	.w5(32'hb9c4a943),
	.w6(32'hbc5bd732),
	.w7(32'hbb8ad604),
	.w8(32'hbc0630a9),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca6b5a8),
	.w1(32'hbc774e9a),
	.w2(32'hbc8b8ab2),
	.w3(32'hbc87d20e),
	.w4(32'hbbba27e0),
	.w5(32'h3b89bc56),
	.w6(32'hbcc2bde4),
	.w7(32'h38116538),
	.w8(32'hbb834c75),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa1e64d),
	.w1(32'hbb4efac8),
	.w2(32'hbad5a90c),
	.w3(32'h3bd96325),
	.w4(32'h3bb5721f),
	.w5(32'h39a3634e),
	.w6(32'hbb358d47),
	.w7(32'hbbb5f3a5),
	.w8(32'hbbb4ff1c),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b09a929),
	.w1(32'h3bd40720),
	.w2(32'hb9235f24),
	.w3(32'hbb124b09),
	.w4(32'h3b2dd35f),
	.w5(32'h3bc9c347),
	.w6(32'hbb986d80),
	.w7(32'h3ba95288),
	.w8(32'hb9050d0f),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbc16b3),
	.w1(32'hbba58881),
	.w2(32'hbbe584ee),
	.w3(32'hbb790151),
	.w4(32'hbb1e884c),
	.w5(32'hbb93b1dc),
	.w6(32'hbbc23a60),
	.w7(32'hbc017407),
	.w8(32'hbb8ae3a3),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd4d00b),
	.w1(32'h3b22c490),
	.w2(32'h3be4ce1a),
	.w3(32'hbbc59142),
	.w4(32'h3b27fd83),
	.w5(32'h3b9613bf),
	.w6(32'hbb90ec18),
	.w7(32'h39a0f059),
	.w8(32'h3b012f91),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6215c2),
	.w1(32'hbc553364),
	.w2(32'hbbf8a0b5),
	.w3(32'h3b4740ed),
	.w4(32'hbbf454f2),
	.w5(32'hbc3932c3),
	.w6(32'h3b4e99da),
	.w7(32'hbb24df3f),
	.w8(32'h395e3716),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc03ed71),
	.w1(32'h3a35c052),
	.w2(32'hbb780329),
	.w3(32'hbbc78fc8),
	.w4(32'h3bca604e),
	.w5(32'h3be53e9d),
	.w6(32'hbbb12227),
	.w7(32'hba3fc458),
	.w8(32'hb9ca0b53),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb2c9ea),
	.w1(32'h39c77904),
	.w2(32'h3aa0f4c5),
	.w3(32'h3bdcd548),
	.w4(32'h3b095939),
	.w5(32'h3bea524e),
	.w6(32'h3ae46f62),
	.w7(32'h3b444c01),
	.w8(32'h3b1d40e6),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0e80a1),
	.w1(32'h3906d040),
	.w2(32'hbb26c5e3),
	.w3(32'h3ab7a9c5),
	.w4(32'h3a6ce27f),
	.w5(32'hbb280b4f),
	.w6(32'hbbb52e8c),
	.w7(32'hbbceadbf),
	.w8(32'hbbb98c3b),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a75230b),
	.w1(32'h397661d5),
	.w2(32'hbbce3ae3),
	.w3(32'hbb777192),
	.w4(32'h3bbad24d),
	.w5(32'hbc11f9e5),
	.w6(32'hbb094e61),
	.w7(32'hbb70b411),
	.w8(32'hbc81ef20),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b81610b),
	.w1(32'hbaabb6a4),
	.w2(32'hbc0212d7),
	.w3(32'h3aaa324d),
	.w4(32'hbb91f90a),
	.w5(32'hbc5e866a),
	.w6(32'h3b02ac84),
	.w7(32'hbb8d7066),
	.w8(32'hbc0feb81),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0dd09b),
	.w1(32'h3b958a08),
	.w2(32'h39b9323c),
	.w3(32'hbbd2456d),
	.w4(32'hbaa795d3),
	.w5(32'h3affce0c),
	.w6(32'hba9030aa),
	.w7(32'hba6c7662),
	.w8(32'h3aedc32f),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4dcd55),
	.w1(32'hbb940236),
	.w2(32'h3ac44b02),
	.w3(32'h3bf4d29f),
	.w4(32'hbbc4a8bc),
	.w5(32'h3bd08c62),
	.w6(32'h3a393ad6),
	.w7(32'hbb0a528d),
	.w8(32'hb9739140),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1173ba),
	.w1(32'hbb172c6b),
	.w2(32'hbb4d1a61),
	.w3(32'h3b267160),
	.w4(32'hbb3c5286),
	.w5(32'hbbba6817),
	.w6(32'hba5b1c5f),
	.w7(32'hbbc090ee),
	.w8(32'hbbd6ff1c),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b01e192),
	.w1(32'hbbc20859),
	.w2(32'hbc5b30d5),
	.w3(32'h3b3cf5af),
	.w4(32'h3b23dd26),
	.w5(32'hbc0328d8),
	.w6(32'hbc2e9dea),
	.w7(32'hbb82727c),
	.w8(32'hbc651034),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5e9b15),
	.w1(32'hbb8097a0),
	.w2(32'hbc2f21e4),
	.w3(32'h3870b11e),
	.w4(32'h3bc8e563),
	.w5(32'hbbac052b),
	.w6(32'h3bcabf20),
	.w7(32'h391ddcc5),
	.w8(32'hbc71a45e),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba73a1e),
	.w1(32'hbbcda437),
	.w2(32'h3afb4fab),
	.w3(32'hbb880080),
	.w4(32'hbbb5e197),
	.w5(32'h3bcc4f98),
	.w6(32'hbbc4def7),
	.w7(32'hbbba0644),
	.w8(32'hb986b17a),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbac634a),
	.w1(32'hb9feb1a4),
	.w2(32'h3b4cdab2),
	.w3(32'h39e32891),
	.w4(32'hbacd0fe9),
	.w5(32'hbaf1eb37),
	.w6(32'hbb3df544),
	.w7(32'hbbc8c36c),
	.w8(32'hbbfc2a56),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7e8d83),
	.w1(32'hb9e6a352),
	.w2(32'h3bddce38),
	.w3(32'h3b5a8008),
	.w4(32'hbb0e3760),
	.w5(32'h3c6b8482),
	.w6(32'hbb4b2ae4),
	.w7(32'hbbf473ae),
	.w8(32'hbb347859),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4c275d),
	.w1(32'hbb8cb873),
	.w2(32'hbb9e3952),
	.w3(32'h3bee87ff),
	.w4(32'h3aefccea),
	.w5(32'hbaa8cb06),
	.w6(32'hbbb4898c),
	.w7(32'hbabbb1f9),
	.w8(32'hbbb3ffc5),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0f46f6),
	.w1(32'hbc5b09cd),
	.w2(32'hbc90e7e5),
	.w3(32'hbc07a63d),
	.w4(32'hbbaf2371),
	.w5(32'hbc22b518),
	.w6(32'hbc0dcbfa),
	.w7(32'hbc31af87),
	.w8(32'hbc63fbb9),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc430490),
	.w1(32'hbc57bf9f),
	.w2(32'hbcb536de),
	.w3(32'h3b8504a1),
	.w4(32'h3abad78f),
	.w5(32'hbc073735),
	.w6(32'hbb4bbf1b),
	.w7(32'hbb0c3cb2),
	.w8(32'hbc662d36),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbad126b),
	.w1(32'h39ebb1c6),
	.w2(32'h392becbf),
	.w3(32'hba8c7bd0),
	.w4(32'h3bb875f6),
	.w5(32'h3bb2377c),
	.w6(32'h3aeec079),
	.w7(32'hba0bcd98),
	.w8(32'hb93d9ed2),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4d3e21),
	.w1(32'hbbdc4202),
	.w2(32'hbbab9e11),
	.w3(32'hba6bebec),
	.w4(32'h3950a73e),
	.w5(32'h3b4b23e3),
	.w6(32'hbb9cace8),
	.w7(32'hbb816b64),
	.w8(32'hbc0075f7),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8f144c),
	.w1(32'hbc1d6d35),
	.w2(32'hbc09e93b),
	.w3(32'h3a1182f9),
	.w4(32'hbb504bd2),
	.w5(32'h3b7b1bf2),
	.w6(32'hbbb4ea09),
	.w7(32'h3623c3be),
	.w8(32'hbc4ab931),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5684ef),
	.w1(32'h3bdc142f),
	.w2(32'h3c1d6535),
	.w3(32'hbb897022),
	.w4(32'h3b94f4cf),
	.w5(32'h3be1e9ee),
	.w6(32'hbc97a0aa),
	.w7(32'hbc14e757),
	.w8(32'hbb81590b),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaa941c),
	.w1(32'hbb8203df),
	.w2(32'hbbd2760f),
	.w3(32'h39851b39),
	.w4(32'hbb45aa61),
	.w5(32'hbbc4d28b),
	.w6(32'hbc0e068b),
	.w7(32'hbb426e62),
	.w8(32'hbc0e6d54),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac08597),
	.w1(32'hbbec7fe3),
	.w2(32'hbb9811a8),
	.w3(32'hb957a570),
	.w4(32'hbc4791e8),
	.w5(32'h3c2b6e4f),
	.w6(32'hb99b040e),
	.w7(32'hbc120473),
	.w8(32'hbbd85b25),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9c274a),
	.w1(32'h3c074b51),
	.w2(32'h3b506404),
	.w3(32'h3caaeda7),
	.w4(32'h3b869a42),
	.w5(32'hbc1a2ee9),
	.w6(32'h3c3da9ad),
	.w7(32'hbbe04149),
	.w8(32'hbc833868),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0f52e9),
	.w1(32'h3ad6dffc),
	.w2(32'hbbaf79fb),
	.w3(32'hbbdee2b4),
	.w4(32'h3bc17e54),
	.w5(32'hbb34d189),
	.w6(32'hbbc404cc),
	.w7(32'h3abf8fdc),
	.w8(32'hbb9404d3),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf9f66b),
	.w1(32'h3b596f07),
	.w2(32'hbb1e398a),
	.w3(32'h3b85c850),
	.w4(32'h3b63d413),
	.w5(32'h3b4db4dc),
	.w6(32'h3aaa82b5),
	.w7(32'hba1e5a29),
	.w8(32'h3af842a8),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbd492a),
	.w1(32'h396f7110),
	.w2(32'hbae2064a),
	.w3(32'hbbbd9112),
	.w4(32'hba2e7413),
	.w5(32'h3a155a96),
	.w6(32'hbb8a033a),
	.w7(32'h3bc7028b),
	.w8(32'h3b03b33d),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc52e8ad),
	.w1(32'hbb7524bf),
	.w2(32'hbb2cc2b4),
	.w3(32'hbaf5e759),
	.w4(32'h3bbb866f),
	.w5(32'h3b07f5bd),
	.w6(32'hbb70c325),
	.w7(32'h3a47a467),
	.w8(32'hbb993ca5),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc23d214),
	.w1(32'h3b1635b5),
	.w2(32'hb9bae56b),
	.w3(32'hbbdc3d11),
	.w4(32'h3bae0dfd),
	.w5(32'h3b608522),
	.w6(32'hbc230db5),
	.w7(32'hbbb2a247),
	.w8(32'hbbbaaa36),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb30c067),
	.w1(32'hbbca2843),
	.w2(32'hbc99fc9d),
	.w3(32'h3bd3de54),
	.w4(32'h39085daa),
	.w5(32'hbc77463c),
	.w6(32'hba98bce3),
	.w7(32'h3a83f6d5),
	.w8(32'hbc923cd7),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc4c297),
	.w1(32'h3ab58e15),
	.w2(32'h3b302d56),
	.w3(32'hbbdab322),
	.w4(32'h3b7f4ae7),
	.w5(32'hbae376c1),
	.w6(32'hbc1fc3d2),
	.w7(32'h3b2a178b),
	.w8(32'h3b8ff283),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd831df),
	.w1(32'hbc5e1a2a),
	.w2(32'hbcac693d),
	.w3(32'h3b986ba0),
	.w4(32'hbb835112),
	.w5(32'hbc785e6f),
	.w6(32'h3ba50846),
	.w7(32'hbc1dfc39),
	.w8(32'hbc8ee2ee),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3fd179),
	.w1(32'h3905fada),
	.w2(32'hbba64661),
	.w3(32'hba010452),
	.w4(32'hbb289170),
	.w5(32'hbb8f8d5e),
	.w6(32'hbb7d3f7c),
	.w7(32'hbbff36cd),
	.w8(32'hbc234bff),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8ad580),
	.w1(32'hbc1cdf1c),
	.w2(32'hbbda6952),
	.w3(32'hbb9542aa),
	.w4(32'hbb08e44f),
	.w5(32'h3c203a1a),
	.w6(32'hbc1398d4),
	.w7(32'h39a3df3a),
	.w8(32'hbaca5f74),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1e60da),
	.w1(32'hbc172805),
	.w2(32'hbc1bb7ca),
	.w3(32'h3bf64b57),
	.w4(32'hbb7606ab),
	.w5(32'hbc5b0c7c),
	.w6(32'h3c4e9965),
	.w7(32'hbc8209da),
	.w8(32'hbcc53a3d),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9f5a44),
	.w1(32'hbb512b5e),
	.w2(32'hbc398efe),
	.w3(32'hbc0ffff6),
	.w4(32'hba7cedf0),
	.w5(32'hbc213513),
	.w6(32'hbc36aba9),
	.w7(32'hbbede444),
	.w8(32'hbc2dec1b),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab51538),
	.w1(32'h3b87c614),
	.w2(32'hbb1b6b63),
	.w3(32'hbaa58405),
	.w4(32'h3b82b2dc),
	.w5(32'hbb5a64bf),
	.w6(32'hbbeaefb8),
	.w7(32'hb92f1b0a),
	.w8(32'h392c6e21),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc05274b),
	.w1(32'h3b152b41),
	.w2(32'h3ada0f09),
	.w3(32'hb9a2c053),
	.w4(32'h39a3479c),
	.w5(32'h3b0549a4),
	.w6(32'h3b57b363),
	.w7(32'hbb9e7e6d),
	.w8(32'hbb7eb15c),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbba70d0),
	.w1(32'hbb79dc95),
	.w2(32'hbc541376),
	.w3(32'hbb8f3c26),
	.w4(32'hbade3c78),
	.w5(32'hbc1ce8da),
	.w6(32'hbc0a4975),
	.w7(32'hbbab4ab4),
	.w8(32'hbc231c6d),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfa3ac2),
	.w1(32'h3be29ed1),
	.w2(32'h3bbf624a),
	.w3(32'hbb5c1f70),
	.w4(32'h3be77906),
	.w5(32'h3947965c),
	.w6(32'h3abc1def),
	.w7(32'h3b10cd35),
	.w8(32'h3b102e2f),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6b21ec),
	.w1(32'hbb2e1a9c),
	.w2(32'hba8de0c8),
	.w3(32'h3b7def9e),
	.w4(32'h3c10370b),
	.w5(32'h3be6a00c),
	.w6(32'h3bcd9c9c),
	.w7(32'h3b9d304a),
	.w8(32'hbaff62eb),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb69b46e),
	.w1(32'h38aa391f),
	.w2(32'h3a98bb64),
	.w3(32'hba1d3e06),
	.w4(32'h3b1f2dc0),
	.w5(32'h3c115bb1),
	.w6(32'hbb6d0661),
	.w7(32'hbabfd35c),
	.w8(32'hbae26e14),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3a2d1f),
	.w1(32'hbb87b631),
	.w2(32'hbb5b1286),
	.w3(32'h3b2dbdc2),
	.w4(32'hb9b10e07),
	.w5(32'h3ae6d32c),
	.w6(32'hbbdd34a2),
	.w7(32'hbbe7fca6),
	.w8(32'hbc805b55),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e53475),
	.w1(32'hbb604ac1),
	.w2(32'hbb87f667),
	.w3(32'hbb796a47),
	.w4(32'hbb14025e),
	.w5(32'hbbfc2666),
	.w6(32'hbb6a3d47),
	.w7(32'hbaef0e66),
	.w8(32'hbbe93cac),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b47d699),
	.w1(32'hb99eddb3),
	.w2(32'h3a8b96fd),
	.w3(32'hbbe913ab),
	.w4(32'h3b9d7d6c),
	.w5(32'h3a294a7f),
	.w6(32'hbc2238a5),
	.w7(32'h3a81e755),
	.w8(32'hba820de2),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba032c6a),
	.w1(32'h3b29dc0d),
	.w2(32'h3ba83240),
	.w3(32'hbb8a024a),
	.w4(32'h3b5dd5b5),
	.w5(32'h3be918c8),
	.w6(32'hbb25de22),
	.w7(32'h3a270eae),
	.w8(32'h3b79d23d),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba3ec4c),
	.w1(32'hbb2f7d9c),
	.w2(32'h3ab10aa0),
	.w3(32'h3c3c2868),
	.w4(32'hbbf60731),
	.w5(32'hbb68ded1),
	.w6(32'h3b6c0b6d),
	.w7(32'hbb74920c),
	.w8(32'hbb680c21),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c43f712),
	.w1(32'h3b0ff711),
	.w2(32'h3c2299e6),
	.w3(32'h3c562815),
	.w4(32'h3aec6330),
	.w5(32'h3c9f7bdd),
	.w6(32'h3c8114bf),
	.w7(32'h3891535e),
	.w8(32'h3c1422ff),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba861ac6),
	.w1(32'hbba39801),
	.w2(32'hbbbab450),
	.w3(32'h3b875e66),
	.w4(32'hbabdadf6),
	.w5(32'hbb9ec45c),
	.w6(32'h3aff5945),
	.w7(32'hba5d2f0e),
	.w8(32'hbba9187c),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabd8730),
	.w1(32'h3a9bd402),
	.w2(32'hba1fb18a),
	.w3(32'hbb9e2919),
	.w4(32'h3b150448),
	.w5(32'h3c0886be),
	.w6(32'hbba719dc),
	.w7(32'hbb185bb2),
	.w8(32'h3a99ff67),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae193cb),
	.w1(32'h3bc362f0),
	.w2(32'hbc057533),
	.w3(32'h3ade8392),
	.w4(32'h3c4f97b8),
	.w5(32'hbc12571b),
	.w6(32'hbcb4a262),
	.w7(32'h3c0fa6cf),
	.w8(32'hbc11f8f1),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a77ce95),
	.w1(32'hbb6d2377),
	.w2(32'hbb71f29e),
	.w3(32'hb8e9c04d),
	.w4(32'hbb724fca),
	.w5(32'hbb55440d),
	.w6(32'h3b08df2e),
	.w7(32'hbb825e03),
	.w8(32'hbb15ebca),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd8a37f),
	.w1(32'h3b9f9ec5),
	.w2(32'h3b689245),
	.w3(32'h3ae92f59),
	.w4(32'h3a84ddb6),
	.w5(32'h3c891300),
	.w6(32'h3c0621a6),
	.w7(32'hbb9f9dcc),
	.w8(32'hbb979c55),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb925acbe),
	.w1(32'hbb2ac62c),
	.w2(32'hbb91a95b),
	.w3(32'h3b97cf00),
	.w4(32'h39745501),
	.w5(32'hbb0ed990),
	.w6(32'h3b279356),
	.w7(32'hba0f9b49),
	.w8(32'h38829832),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc557a42),
	.w1(32'hbb9af1f0),
	.w2(32'hbc544fa3),
	.w3(32'hbb5b5700),
	.w4(32'h3c0bbbfd),
	.w5(32'h3b584b43),
	.w6(32'hbc039198),
	.w7(32'h3b6cb70e),
	.w8(32'hbc14016d),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe44d0e),
	.w1(32'h3ab519f4),
	.w2(32'hbc042e7e),
	.w3(32'hbb5bccbe),
	.w4(32'h3be2f9d6),
	.w5(32'h3acd95da),
	.w6(32'hbbf5e89a),
	.w7(32'h3a0a5734),
	.w8(32'hbbbf1f12),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0fd951),
	.w1(32'hbc272d82),
	.w2(32'hbcb711a5),
	.w3(32'hbc48a721),
	.w4(32'hbbe629e7),
	.w5(32'hbc9a150c),
	.w6(32'hbc1c9053),
	.w7(32'hbbeb1459),
	.w8(32'hbc974f9a),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3913701a),
	.w1(32'h3b45768a),
	.w2(32'hba8df3a0),
	.w3(32'hbb924296),
	.w4(32'h3b9af9fa),
	.w5(32'hb9a4571a),
	.w6(32'hbb09b8c4),
	.w7(32'h3b90efcc),
	.w8(32'h3ae2b332),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb87df0),
	.w1(32'hbc0a48b7),
	.w2(32'hbc1f491e),
	.w3(32'hbb550f73),
	.w4(32'h3b6097e1),
	.w5(32'hbbb9a206),
	.w6(32'hbaea0fdd),
	.w7(32'hbab7f368),
	.w8(32'hbba5908e),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b377d89),
	.w1(32'hbb24546c),
	.w2(32'hbb57f258),
	.w3(32'h3a106b3e),
	.w4(32'hbaa133eb),
	.w5(32'hba6ed7b4),
	.w6(32'h3a535ef6),
	.w7(32'hbbbb2102),
	.w8(32'h3b649910),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3c1743),
	.w1(32'h3ab05b08),
	.w2(32'hbbcdbe0c),
	.w3(32'h3c04ac9c),
	.w4(32'h3a62cae4),
	.w5(32'h3b21ef71),
	.w6(32'h398741ec),
	.w7(32'h3a8cc494),
	.w8(32'hbb814669),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba75de1),
	.w1(32'hba26d0c8),
	.w2(32'h3ad9df9a),
	.w3(32'h3b1994bb),
	.w4(32'h3a9b63c4),
	.w5(32'hbbc8bf44),
	.w6(32'hbb27240d),
	.w7(32'h3b7d4567),
	.w8(32'hbb0fa737),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0528fa),
	.w1(32'hbc16f9f0),
	.w2(32'hbc1e7bce),
	.w3(32'hbba1a67a),
	.w4(32'h3a5a5eed),
	.w5(32'hbbbaeb2d),
	.w6(32'hbc222af9),
	.w7(32'hba3d2f66),
	.w8(32'hbc11c0ac),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0f1cff),
	.w1(32'hbaecb19d),
	.w2(32'h3bb2f050),
	.w3(32'hbb1969c5),
	.w4(32'h3b91eb21),
	.w5(32'h3c096e4d),
	.w6(32'hba89fee4),
	.w7(32'h3bd8fd30),
	.w8(32'h3be07508),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b923dc3),
	.w1(32'hbb9e07d0),
	.w2(32'h3aade3cb),
	.w3(32'h3b6e0cde),
	.w4(32'hbb0dd023),
	.w5(32'h3c3d994b),
	.w6(32'h3bcfc397),
	.w7(32'hb9b6fc1c),
	.w8(32'h38aee171),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab6dd00),
	.w1(32'hbb6c420b),
	.w2(32'hbaa55858),
	.w3(32'hbb707ece),
	.w4(32'hbae477ac),
	.w5(32'h3c1e0ff7),
	.w6(32'hbb2496ba),
	.w7(32'hbbd97573),
	.w8(32'hbbdf90d7),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc57f754),
	.w1(32'h3b088128),
	.w2(32'hbbdb8c38),
	.w3(32'hbbf3e8e8),
	.w4(32'h3b9f57b5),
	.w5(32'hbb5f8154),
	.w6(32'hbc3a73d4),
	.w7(32'h3b2f9d45),
	.w8(32'hbc19212e),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6c82a0),
	.w1(32'hbc730800),
	.w2(32'hbbfbd94c),
	.w3(32'hbba2dbab),
	.w4(32'hbc2c2928),
	.w5(32'hbb2f75ae),
	.w6(32'hbb4037f0),
	.w7(32'hbbd1f254),
	.w8(32'hbbba0b2a),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9145ea),
	.w1(32'h3b7337a3),
	.w2(32'hbbb58c96),
	.w3(32'h3af17404),
	.w4(32'h3b12e79b),
	.w5(32'hbb977c54),
	.w6(32'hba55e906),
	.w7(32'h3b851f92),
	.w8(32'hbc1b6961),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc93cddf),
	.w1(32'hbc4eb5a4),
	.w2(32'hbcdb8739),
	.w3(32'hbc0adb3c),
	.w4(32'h3bb60e75),
	.w5(32'hbc42c33c),
	.w6(32'hbc795d94),
	.w7(32'hbbfb0de5),
	.w8(32'hbc94dd8f),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabeb561),
	.w1(32'h3aed55ff),
	.w2(32'hbc640a43),
	.w3(32'hbb9228d3),
	.w4(32'h3c4dbc37),
	.w5(32'h3b34e036),
	.w6(32'hba3d498a),
	.w7(32'hbb31cc32),
	.w8(32'hbc6defb9),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc159f55),
	.w1(32'hbb4f081d),
	.w2(32'hbc23fb84),
	.w3(32'hbb4965e6),
	.w4(32'hbbbb9156),
	.w5(32'hbc1f30d4),
	.w6(32'hbba25138),
	.w7(32'hbba5bda9),
	.w8(32'hbbe0dde9),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaab75a),
	.w1(32'hbb47996a),
	.w2(32'hbac034e7),
	.w3(32'hbbdc02e3),
	.w4(32'hbb13e295),
	.w5(32'h3c27063a),
	.w6(32'hbb8ce900),
	.w7(32'hbb48bae1),
	.w8(32'hbb2bdc8d),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb898b91),
	.w1(32'h3b9001f0),
	.w2(32'hb90e757b),
	.w3(32'hbabf0631),
	.w4(32'h3b2deacc),
	.w5(32'h38c106c9),
	.w6(32'hbbd4cf2c),
	.w7(32'h3ba152b4),
	.w8(32'hbb1861d7),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3fd3d1),
	.w1(32'h3bff655d),
	.w2(32'h3b99b151),
	.w3(32'hbb0c40cc),
	.w4(32'h3bd04744),
	.w5(32'h3b88a9ce),
	.w6(32'hbba66351),
	.w7(32'h3bbf1d56),
	.w8(32'h3b337ce7),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb03bd51),
	.w1(32'hbc18bf46),
	.w2(32'hbc323903),
	.w3(32'hba6f142a),
	.w4(32'hbbd7ebdf),
	.w5(32'hbc5d4963),
	.w6(32'hbbaf2450),
	.w7(32'hbb695664),
	.w8(32'hbc112739),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4fa7ab),
	.w1(32'h3ad99d19),
	.w2(32'hba955b2c),
	.w3(32'hbb96e8eb),
	.w4(32'h3b8fa51a),
	.w5(32'h3acc5c71),
	.w6(32'hbbd50879),
	.w7(32'hbb8ae499),
	.w8(32'hbb834a35),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7ce04f),
	.w1(32'hbbc083f0),
	.w2(32'hbc6c3a6a),
	.w3(32'h3ab550dd),
	.w4(32'hbb0b311a),
	.w5(32'hbbb7bb4f),
	.w6(32'hbaf54f5d),
	.w7(32'hbb8bc732),
	.w8(32'hbc517654),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8932db),
	.w1(32'hbb472742),
	.w2(32'hbb84e74e),
	.w3(32'h3a888341),
	.w4(32'hbb1201fd),
	.w5(32'h3a25044c),
	.w6(32'h3ac4e330),
	.w7(32'hba89128f),
	.w8(32'hba5133b4),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b44bbe8),
	.w1(32'hbb9979c9),
	.w2(32'hbca47afd),
	.w3(32'h3c93e43d),
	.w4(32'h3c515de7),
	.w5(32'hbc20fd1e),
	.w6(32'h3c093419),
	.w7(32'h3b0f226e),
	.w8(32'hbc9fc70a),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5804ab),
	.w1(32'hbb9df239),
	.w2(32'hbb4d08ee),
	.w3(32'hbb60a630),
	.w4(32'h3b2c35b0),
	.w5(32'hbaf20f84),
	.w6(32'hbbd0e1e3),
	.w7(32'h3b7f9bb1),
	.w8(32'h3b0d2083),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3968d415),
	.w1(32'hba7f22fb),
	.w2(32'h3b4a31db),
	.w3(32'h3b246734),
	.w4(32'h3bf8ff10),
	.w5(32'h3b8c5c0e),
	.w6(32'hb97f1702),
	.w7(32'hba0367b1),
	.w8(32'h39bf3661),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba2a804),
	.w1(32'hbc85eca2),
	.w2(32'hbc4406b7),
	.w3(32'h3bbb69c6),
	.w4(32'hbc0ea58a),
	.w5(32'hbbff4819),
	.w6(32'hbb6c8bde),
	.w7(32'hba00d53b),
	.w8(32'h3b9962d4),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb607c8d),
	.w1(32'hbb0fc451),
	.w2(32'h3bc1b741),
	.w3(32'hbc08eba8),
	.w4(32'h3bb9b47a),
	.w5(32'h3c39b0bb),
	.w6(32'hbba1f51b),
	.w7(32'h3b802d58),
	.w8(32'h3b612c25),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7aca24),
	.w1(32'hbb5b1832),
	.w2(32'hbc26bbde),
	.w3(32'h3bafd3fd),
	.w4(32'h3ba86571),
	.w5(32'hbb85cb48),
	.w6(32'h3a50dd42),
	.w7(32'hbad47fc5),
	.w8(32'hbbff5722),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba639473),
	.w1(32'hbbd50d51),
	.w2(32'hbc857f08),
	.w3(32'hbb08a779),
	.w4(32'h39b6a0ca),
	.w5(32'hbc811e7e),
	.w6(32'hbb8ad8c3),
	.w7(32'hbbab2c3e),
	.w8(32'hbc93eb69),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbed9e37),
	.w1(32'hbab6b4af),
	.w2(32'hbc07f67e),
	.w3(32'hbb50509e),
	.w4(32'h3aa2c274),
	.w5(32'h3b033da4),
	.w6(32'hbc4b4611),
	.w7(32'hbc58512d),
	.w8(32'hbc80d0d6),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf0b278),
	.w1(32'h39f7cd1c),
	.w2(32'hbbac76f6),
	.w3(32'hbc3f6f15),
	.w4(32'h3ba93c26),
	.w5(32'h39ab95f9),
	.w6(32'hbbf4d1a8),
	.w7(32'hbb9c6b1b),
	.w8(32'h3baa6d50),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb419e10),
	.w1(32'h3a96ab56),
	.w2(32'hbbfebf7f),
	.w3(32'h3a79f8cc),
	.w4(32'h3c38c0b9),
	.w5(32'h3b219d7b),
	.w6(32'hbbd2b141),
	.w7(32'h3ae58fd1),
	.w8(32'hbc0725a4),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd08f48),
	.w1(32'hbc2a0bd1),
	.w2(32'hbc1772df),
	.w3(32'hbb8f6dc0),
	.w4(32'hbb853984),
	.w5(32'hbb947aca),
	.w6(32'hbb560dc9),
	.w7(32'hbc204179),
	.w8(32'hbc03795d),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc52387b),
	.w1(32'hbc5d6b7a),
	.w2(32'hbccee27a),
	.w3(32'h3b081f2a),
	.w4(32'h3bfb8283),
	.w5(32'h3b218271),
	.w6(32'hbba70894),
	.w7(32'hbb7097b6),
	.w8(32'hbc5eca90),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc55a303),
	.w1(32'hbba2d4ca),
	.w2(32'hbbc46830),
	.w3(32'hbb37dea3),
	.w4(32'hbc141ffe),
	.w5(32'hbbbb8538),
	.w6(32'hbbc00eaa),
	.w7(32'hbb8c8473),
	.w8(32'hbb6f6db0),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba67103),
	.w1(32'hbbb24f26),
	.w2(32'hbbeb2100),
	.w3(32'hbb6b9db3),
	.w4(32'hbb17b885),
	.w5(32'hbb100b78),
	.w6(32'hbbcb702b),
	.w7(32'hbbb87704),
	.w8(32'hbc3576f7),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc9501e),
	.w1(32'hbc7cf8b0),
	.w2(32'hbbd8db61),
	.w3(32'h3b854fcf),
	.w4(32'hb92884ae),
	.w5(32'hbb81a7dc),
	.w6(32'hbca2cecc),
	.w7(32'hbb49e799),
	.w8(32'hbc5ce33d),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadd99bd),
	.w1(32'h3b5b7645),
	.w2(32'hbbce9c89),
	.w3(32'hbb39fa7d),
	.w4(32'h3ba14f62),
	.w5(32'hba7cdb4f),
	.w6(32'hbc8b2c54),
	.w7(32'hbbcbbd94),
	.w8(32'hbc5538c6),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcaefa4),
	.w1(32'h3c7c9355),
	.w2(32'h3b8b7db0),
	.w3(32'hbb67d670),
	.w4(32'h3c32e168),
	.w5(32'hba992d56),
	.w6(32'hbc6a91fd),
	.w7(32'hbaa63449),
	.w8(32'hbc298847),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e41d60),
	.w1(32'hbc5699a3),
	.w2(32'hbc3aec6b),
	.w3(32'h3b835cfb),
	.w4(32'hb8fb504b),
	.w5(32'hbc4b1e4f),
	.w6(32'h3bbfa2ae),
	.w7(32'hbc099ee1),
	.w8(32'hbc40684f),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb705219),
	.w1(32'hbc0c1910),
	.w2(32'hba767d25),
	.w3(32'hbaccde62),
	.w4(32'hbbf4014d),
	.w5(32'hbbfc117d),
	.w6(32'hbc16c307),
	.w7(32'hbc0af883),
	.w8(32'hbc76e67b),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc166b18),
	.w1(32'hbb521cda),
	.w2(32'h3c082701),
	.w3(32'hbb508b3f),
	.w4(32'hba5a4205),
	.w5(32'h3baf1bba),
	.w6(32'hbc3eef6a),
	.w7(32'hbb20e37d),
	.w8(32'hbb9b50e1),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd01976),
	.w1(32'hbba10cd3),
	.w2(32'hbc9f82f5),
	.w3(32'h3b157671),
	.w4(32'hbbad00e3),
	.w5(32'hbc25ad82),
	.w6(32'hbc1c5ddd),
	.w7(32'hbb1d8123),
	.w8(32'hbbacff20),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc393d87),
	.w1(32'h3b35b7e8),
	.w2(32'h3aed1004),
	.w3(32'h3ad13dfe),
	.w4(32'h3b896989),
	.w5(32'h3c9296e1),
	.w6(32'hbc15aca3),
	.w7(32'h3aa30f78),
	.w8(32'hbb341358),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2aa899),
	.w1(32'h3bbad090),
	.w2(32'h3b323ce1),
	.w3(32'h3c734031),
	.w4(32'hba6b344d),
	.w5(32'hbb8ef825),
	.w6(32'hbb36fa01),
	.w7(32'hbaac79df),
	.w8(32'hbc48e1f1),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3c88e5),
	.w1(32'h3c0346c0),
	.w2(32'h3bcf381f),
	.w3(32'hbb14dad1),
	.w4(32'h3c4f6ad7),
	.w5(32'h3c545b71),
	.w6(32'h3a333512),
	.w7(32'h3b1990e5),
	.w8(32'hbba45a61),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39584a36),
	.w1(32'hbb347f0c),
	.w2(32'hba8d2500),
	.w3(32'h3b8c73cd),
	.w4(32'h3ba1bdef),
	.w5(32'h3af655a6),
	.w6(32'hb9fc6717),
	.w7(32'hbb44295a),
	.w8(32'hbc059f2c),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b86a0d4),
	.w1(32'hb9d18926),
	.w2(32'hba6e5ed5),
	.w3(32'h3a6ab6e3),
	.w4(32'h3b7ce1b2),
	.w5(32'hbb9127bd),
	.w6(32'h3be61f77),
	.w7(32'hbbe47aab),
	.w8(32'hbbe6109d),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb022145),
	.w1(32'hb9372d91),
	.w2(32'h3b05a7b2),
	.w3(32'hbb460ea2),
	.w4(32'hbbc8dca6),
	.w5(32'h3ba4d388),
	.w6(32'hbbf625e1),
	.w7(32'hbbd8f70e),
	.w8(32'h3b5250cc),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2871c1),
	.w1(32'hbb2fe5da),
	.w2(32'h3b162932),
	.w3(32'h3c9311cd),
	.w4(32'hba3cb931),
	.w5(32'hbac245f5),
	.w6(32'h3ba88192),
	.w7(32'hbad8199c),
	.w8(32'hbbce3263),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdd4793),
	.w1(32'h3b563ecd),
	.w2(32'hbba36e9f),
	.w3(32'hbc09d4eb),
	.w4(32'hbad8541a),
	.w5(32'hbc0b6a6f),
	.w6(32'hbbb40274),
	.w7(32'h3ada3c39),
	.w8(32'h3a314849),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb174658),
	.w1(32'hbc05318a),
	.w2(32'hbc4770f4),
	.w3(32'hbb10a433),
	.w4(32'hbc1ddaf2),
	.w5(32'hbc66e6a3),
	.w6(32'h3bab9850),
	.w7(32'hbabccff7),
	.w8(32'hbbb9dbc3),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4ff5be),
	.w1(32'hbc5dd956),
	.w2(32'hbc17b1a4),
	.w3(32'hbc115bad),
	.w4(32'h3b4cb17d),
	.w5(32'h3ad139f6),
	.w6(32'hbc807337),
	.w7(32'hbc72655c),
	.w8(32'hbc5bbfe6),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb90bf5c),
	.w1(32'h3ac68b9a),
	.w2(32'h3bd6ed97),
	.w3(32'h3b13c577),
	.w4(32'h3c614a6e),
	.w5(32'h3c67cef3),
	.w6(32'hbc171b2a),
	.w7(32'h3b56c1c3),
	.w8(32'hbb5e47e1),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b68842b),
	.w1(32'hbb49f562),
	.w2(32'hba82f361),
	.w3(32'h3c1e1bcf),
	.w4(32'h3b01592a),
	.w5(32'h3b37b36a),
	.w6(32'h3b998f00),
	.w7(32'h3a2bd44d),
	.w8(32'hbabb7049),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9b79f5),
	.w1(32'hbc3da8a7),
	.w2(32'hbc23e573),
	.w3(32'hbb364aa6),
	.w4(32'h3c698ae9),
	.w5(32'h3c8aa9cf),
	.w6(32'hbc84928e),
	.w7(32'h3bd78ce4),
	.w8(32'hbabfc096),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a505a3d),
	.w1(32'hb9a82949),
	.w2(32'hbc123928),
	.w3(32'h3c903582),
	.w4(32'h3c2c8866),
	.w5(32'h3bb19d5c),
	.w6(32'hbb37e426),
	.w7(32'h3a5b82a4),
	.w8(32'hbb49aa74),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7352b0),
	.w1(32'hbc083c21),
	.w2(32'hbbed00b3),
	.w3(32'h3b8aa8b2),
	.w4(32'hbb320679),
	.w5(32'hbc258712),
	.w6(32'h3b13edec),
	.w7(32'hbc52e6da),
	.w8(32'hbc93b336),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd8fed2),
	.w1(32'hbbbc76f4),
	.w2(32'hbc2491bf),
	.w3(32'hbb8f062c),
	.w4(32'hbb54e898),
	.w5(32'hbbaae853),
	.w6(32'hbc7f82af),
	.w7(32'hbbfbc59b),
	.w8(32'hbc6bf698),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9726af),
	.w1(32'hbbf17d23),
	.w2(32'hbb517221),
	.w3(32'hbb9e063a),
	.w4(32'hbc001ec4),
	.w5(32'h39bb1940),
	.w6(32'hbbe9d748),
	.w7(32'h3ab53459),
	.w8(32'h3bbee8eb),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8cddff),
	.w1(32'h3bc9de50),
	.w2(32'hbb00013b),
	.w3(32'hbb2c602b),
	.w4(32'h3ba61cf4),
	.w5(32'h3b82a7d2),
	.w6(32'hbbf60be2),
	.w7(32'h3af054e8),
	.w8(32'hb92462ab),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdac3d4),
	.w1(32'hbbf2a433),
	.w2(32'hbb4f8ffe),
	.w3(32'h3ac484b9),
	.w4(32'hbb4c5cb1),
	.w5(32'hbbc699c7),
	.w6(32'h3aad27ff),
	.w7(32'hbbdd0c30),
	.w8(32'hbbd600d0),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac57172),
	.w1(32'h39ae808a),
	.w2(32'hba2d1fc8),
	.w3(32'hbada3916),
	.w4(32'h3b2edb4c),
	.w5(32'h3afa11fb),
	.w6(32'hbc07bbab),
	.w7(32'hbc0b7635),
	.w8(32'hbc386198),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bffc77f),
	.w1(32'h3b6e0e05),
	.w2(32'hbb8077a3),
	.w3(32'h3beef2f7),
	.w4(32'hbba99b41),
	.w5(32'hbac321ac),
	.w6(32'hbb67cd9d),
	.w7(32'h3a414f28),
	.w8(32'hbb412c15),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc77d81d),
	.w1(32'hbc647f22),
	.w2(32'hbcf11765),
	.w3(32'hbbdb27b7),
	.w4(32'h3b4bffac),
	.w5(32'hbc895cde),
	.w6(32'hbc38957e),
	.w7(32'hbbd716ca),
	.w8(32'hbcb78690),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1579b2),
	.w1(32'hbc4542db),
	.w2(32'hbc426cce),
	.w3(32'hbada7b16),
	.w4(32'hba4b4398),
	.w5(32'h3a59aa41),
	.w6(32'hbbc8b8dc),
	.w7(32'hbac1b473),
	.w8(32'hbc03275c),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc82b7cd),
	.w1(32'hbc43e182),
	.w2(32'hbc2994e3),
	.w3(32'hbb3e625d),
	.w4(32'hbb0bc316),
	.w5(32'h3bbca774),
	.w6(32'hbbc5caf5),
	.w7(32'hbc08a6cc),
	.w8(32'hbc205fc9),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba114dba),
	.w1(32'h3bf04534),
	.w2(32'h3bb5dffc),
	.w3(32'h36f7a1ec),
	.w4(32'h3bc429ac),
	.w5(32'h3c439c8f),
	.w6(32'hbb503d72),
	.w7(32'h3b74f9d2),
	.w8(32'hb8f9bcf7),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae25dfc),
	.w1(32'hbbe74965),
	.w2(32'hbc213963),
	.w3(32'hbafd4e1e),
	.w4(32'hbbcaae18),
	.w5(32'hbbe060d4),
	.w6(32'hbb5c80b6),
	.w7(32'hbc03431b),
	.w8(32'hbbbc7917),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc05092f),
	.w1(32'hbbb905ff),
	.w2(32'hbb1f2a32),
	.w3(32'hba908c98),
	.w4(32'hbbe5a56b),
	.w5(32'h3ba39cb8),
	.w6(32'hbb426018),
	.w7(32'hbbbd5b51),
	.w8(32'hbb32af24),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc44b202),
	.w1(32'hbae52e9a),
	.w2(32'h3b922040),
	.w3(32'hbc38e7f3),
	.w4(32'h3a1c970c),
	.w5(32'h3be5be06),
	.w6(32'hbc036708),
	.w7(32'h3a6d08d5),
	.w8(32'hbb27b4cf),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc77b236),
	.w1(32'hbc0c17f0),
	.w2(32'hbc06ea68),
	.w3(32'hbad98d49),
	.w4(32'h3be3615a),
	.w5(32'h3b8b69a3),
	.w6(32'hbc074196),
	.w7(32'hbb69367a),
	.w8(32'hbc85dece),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba73e11b),
	.w1(32'h3b6c2bfe),
	.w2(32'h3c714a5c),
	.w3(32'h3b296e31),
	.w4(32'h3b8f3d2d),
	.w5(32'h3c59a453),
	.w6(32'hbbb2e8fc),
	.w7(32'h3bc5487d),
	.w8(32'h3c568979),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c18cb5a),
	.w1(32'h3bb5ab9a),
	.w2(32'h3c09357a),
	.w3(32'h3c21a70a),
	.w4(32'h3b685f42),
	.w5(32'h3bd9d49f),
	.w6(32'h3b9cf7ce),
	.w7(32'h3b2d8b68),
	.w8(32'h3bbec2cb),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae023d1),
	.w1(32'h3bb527aa),
	.w2(32'hba20a425),
	.w3(32'hbbdb90df),
	.w4(32'h3b9806d6),
	.w5(32'hbc03ec06),
	.w6(32'hbad8faa3),
	.w7(32'h3bacc7c1),
	.w8(32'hbc09465b),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aab2982),
	.w1(32'hbc461f40),
	.w2(32'hbbbc9a22),
	.w3(32'h3aeb6394),
	.w4(32'hbc40e3c8),
	.w5(32'hbc66b3f5),
	.w6(32'h3acc8321),
	.w7(32'hbc0e7c39),
	.w8(32'hbc3f299a),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf17dfc),
	.w1(32'hbb51f5da),
	.w2(32'hbc1f6402),
	.w3(32'hbb50c6ed),
	.w4(32'h3be40e8f),
	.w5(32'hba1cca90),
	.w6(32'hbc241d9b),
	.w7(32'h3b2a8632),
	.w8(32'hbbe59e74),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3df516),
	.w1(32'hbc30b327),
	.w2(32'hbc5fab81),
	.w3(32'h3ba3836f),
	.w4(32'hbb2b5bb2),
	.w5(32'hbc7b27df),
	.w6(32'h3a984c8e),
	.w7(32'hbc2ca318),
	.w8(32'hbc91b1e9),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf4edf8),
	.w1(32'hbca00916),
	.w2(32'hbc8fab9d),
	.w3(32'hbc85f4bc),
	.w4(32'h3ae5085c),
	.w5(32'h3c035991),
	.w6(32'hbcef3648),
	.w7(32'hbb0e03e0),
	.w8(32'hbc4a2d47),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac8f0ad),
	.w1(32'h3bdbed45),
	.w2(32'h3ca564e4),
	.w3(32'h3a3b8748),
	.w4(32'h3cc66961),
	.w5(32'h3d261158),
	.w6(32'hbba44293),
	.w7(32'h3bb6b7d8),
	.w8(32'h3c997333),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c77b73d),
	.w1(32'hbb03b314),
	.w2(32'h3c137ade),
	.w3(32'h3caefa77),
	.w4(32'h3b5723dc),
	.w5(32'h3af92895),
	.w6(32'hb99f456c),
	.w7(32'hbbe97956),
	.w8(32'hbc0f6f80),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule