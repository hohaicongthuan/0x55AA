module layer_10_featuremap_124(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88121df),
	.w1(32'h3921c067),
	.w2(32'hb93ec821),
	.w3(32'hb99ac99d),
	.w4(32'h3b1fb494),
	.w5(32'h3a5973a3),
	.w6(32'hb51312fd),
	.w7(32'hb86a49ba),
	.w8(32'h3a1d7cca),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae38737),
	.w1(32'h39ee3085),
	.w2(32'h399950a5),
	.w3(32'hbaa0108a),
	.w4(32'hb9675e32),
	.w5(32'hb9c1f0b3),
	.w6(32'hb8a04c53),
	.w7(32'h38d1c828),
	.w8(32'hba848413),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3677b6fb),
	.w1(32'hb837ef31),
	.w2(32'h3a5afc40),
	.w3(32'hba02805f),
	.w4(32'hb9303d2b),
	.w5(32'h3a28d6ed),
	.w6(32'hb9f9e16f),
	.w7(32'h3944981a),
	.w8(32'hba4ec9c5),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e25ef2),
	.w1(32'hb9de995c),
	.w2(32'h3aaad209),
	.w3(32'hb8d0b7de),
	.w4(32'hba95096b),
	.w5(32'h394a45e4),
	.w6(32'h39ef2b61),
	.w7(32'h39ed438e),
	.w8(32'hba4d67fb),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a4b79e),
	.w1(32'h3a9a8b4c),
	.w2(32'hb9538141),
	.w3(32'hba19e8b8),
	.w4(32'h3aab785e),
	.w5(32'h39abb2b3),
	.w6(32'h3a670ab9),
	.w7(32'h39b635bf),
	.w8(32'h3ad5279b),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac37837),
	.w1(32'hba8c593a),
	.w2(32'hb64145da),
	.w3(32'h3a6352fe),
	.w4(32'hbab5f6df),
	.w5(32'hbaad1628),
	.w6(32'hba60f675),
	.w7(32'hb9faf131),
	.w8(32'hba948216),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba182ade),
	.w1(32'h3aaa6b76),
	.w2(32'h3af4bd53),
	.w3(32'hbad492a6),
	.w4(32'h3a822a0c),
	.w5(32'h3aca9ad5),
	.w6(32'h3a529985),
	.w7(32'h3a9782bd),
	.w8(32'h3a0ee31b),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab8e802),
	.w1(32'h3ae2a7b6),
	.w2(32'h3a9f704e),
	.w3(32'hba47e71e),
	.w4(32'hb80a4fd6),
	.w5(32'hb9fba604),
	.w6(32'hba395907),
	.w7(32'hb941d4e9),
	.w8(32'h39317372),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392c13fd),
	.w1(32'hba35779f),
	.w2(32'hb8cb0613),
	.w3(32'hba8cd065),
	.w4(32'hba8c87f4),
	.w5(32'hba1a1e74),
	.w6(32'hbb0434b4),
	.w7(32'hbac704ea),
	.w8(32'hba3a2578),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0b8c1e),
	.w1(32'h3a5f4a31),
	.w2(32'h3b19a335),
	.w3(32'h39d9f00d),
	.w4(32'h3988240d),
	.w5(32'h3aff42d4),
	.w6(32'hb7cdb941),
	.w7(32'hbab04faa),
	.w8(32'hbac762e0),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3c11c0),
	.w1(32'h395da812),
	.w2(32'h3a83ebd1),
	.w3(32'hba15b16b),
	.w4(32'hbb281fb9),
	.w5(32'hbb69b251),
	.w6(32'hba4680f3),
	.w7(32'h39104156),
	.w8(32'hba1ebf26),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5c7ca9),
	.w1(32'hba7a51ee),
	.w2(32'h39805e48),
	.w3(32'hbbb3a0e7),
	.w4(32'hba6f8dd3),
	.w5(32'hb96d4648),
	.w6(32'hb9b57e48),
	.w7(32'h3aa9154e),
	.w8(32'hb9c451a9),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4323d3),
	.w1(32'h3979ea72),
	.w2(32'h3a55b856),
	.w3(32'hba92e7a4),
	.w4(32'hba38ee17),
	.w5(32'h39905598),
	.w6(32'hba3a9f70),
	.w7(32'hbb08a29d),
	.w8(32'hba546940),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cd474c),
	.w1(32'h3acdaf78),
	.w2(32'h3aaa66f3),
	.w3(32'h391a8191),
	.w4(32'h3ad35376),
	.w5(32'h3a174dae),
	.w6(32'h3afa69e8),
	.w7(32'h3ad5947f),
	.w8(32'h3a373a69),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9f5c0f),
	.w1(32'hbadaabd8),
	.w2(32'hbb18a273),
	.w3(32'hba32d658),
	.w4(32'hbb243a8c),
	.w5(32'hbb04fece),
	.w6(32'h39f8050c),
	.w7(32'hba4a2a85),
	.w8(32'hb9efac28),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38754db5),
	.w1(32'hb884072e),
	.w2(32'h3a08fcb3),
	.w3(32'hba03fc5b),
	.w4(32'hb9d8e0c5),
	.w5(32'h3a18fba1),
	.w6(32'hbab30a9d),
	.w7(32'hbac8f7ec),
	.w8(32'hb8e9fe5a),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91092af),
	.w1(32'hba4f8942),
	.w2(32'h3b258fe5),
	.w3(32'h36e78545),
	.w4(32'h3af19afa),
	.w5(32'h3ba8ab5a),
	.w6(32'hba904896),
	.w7(32'h3b471a65),
	.w8(32'hba875471),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a46fd82),
	.w1(32'h3a9056d8),
	.w2(32'h3b286443),
	.w3(32'h38afab08),
	.w4(32'hba002873),
	.w5(32'h3a896847),
	.w6(32'hba09f836),
	.w7(32'hba3925a6),
	.w8(32'hba010bbb),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39de64f3),
	.w1(32'h3a0b55f9),
	.w2(32'h3ac046e9),
	.w3(32'hba9b22de),
	.w4(32'hb92f161c),
	.w5(32'h3a84b5f9),
	.w6(32'hba76c8a6),
	.w7(32'hb91750d3),
	.w8(32'hb94894e7),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9da90cf),
	.w1(32'hba9b3b8d),
	.w2(32'hba8f18f9),
	.w3(32'hb4857e40),
	.w4(32'hba317524),
	.w5(32'hba8623f9),
	.w6(32'hbaa1551d),
	.w7(32'hba859ed5),
	.w8(32'hba777802),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba851db9),
	.w1(32'h3b51931e),
	.w2(32'h3baad473),
	.w3(32'hba8a065d),
	.w4(32'h3b2f0cea),
	.w5(32'h3b3be558),
	.w6(32'h3b3c16d2),
	.w7(32'h3b64a30c),
	.w8(32'h3a3dfc4e),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aad9d35),
	.w1(32'hba051dc5),
	.w2(32'hbae8b121),
	.w3(32'h3889cf1a),
	.w4(32'h3a07f2e3),
	.w5(32'h3a05a707),
	.w6(32'hba7a1e87),
	.w7(32'h39a70b1f),
	.w8(32'hbaf6ec80),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab58aa1),
	.w1(32'h3c056a9a),
	.w2(32'h3c21b687),
	.w3(32'hba437ceb),
	.w4(32'h3a76c791),
	.w5(32'h3b9ee4fc),
	.w6(32'h3b961b56),
	.w7(32'h3b84c09b),
	.w8(32'h3a03f94b),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0e467f),
	.w1(32'h3a97d686),
	.w2(32'h3a968c63),
	.w3(32'h3b923edf),
	.w4(32'hb90df4fe),
	.w5(32'h385ab603),
	.w6(32'h3a2b9c54),
	.w7(32'hba971e48),
	.w8(32'hb959658d),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e72713),
	.w1(32'hb9e99918),
	.w2(32'hb8058b06),
	.w3(32'hbab43e6a),
	.w4(32'hba5eebaf),
	.w5(32'hbabfb4a6),
	.w6(32'hba94c750),
	.w7(32'hba1b0a44),
	.w8(32'hbb108087),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37fc9b57),
	.w1(32'hbb218e84),
	.w2(32'hbadaf049),
	.w3(32'h39072f75),
	.w4(32'h39a8ff5d),
	.w5(32'h3ad6dead),
	.w6(32'hbb7aeefb),
	.w7(32'hbb5092a1),
	.w8(32'hbb70ff1d),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf3f82a),
	.w1(32'hbaf4743b),
	.w2(32'hbaea54c1),
	.w3(32'h393e1a48),
	.w4(32'hba9a1225),
	.w5(32'hbad50917),
	.w6(32'hbadf9442),
	.w7(32'hbadd5d5a),
	.w8(32'hbaad4178),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb390820),
	.w1(32'h3a01b465),
	.w2(32'h39371653),
	.w3(32'hbb20823b),
	.w4(32'h3ac7164a),
	.w5(32'h39d8ca01),
	.w6(32'h3a9177e7),
	.w7(32'h3ad21aa6),
	.w8(32'h39967914),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa1cd80),
	.w1(32'h3b517b19),
	.w2(32'h3b9303cf),
	.w3(32'hba30af71),
	.w4(32'h3a7771d7),
	.w5(32'h3ab89a21),
	.w6(32'h3b1a8c27),
	.w7(32'h3b87151c),
	.w8(32'hb98a8990),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b991a43),
	.w1(32'h3ba018ba),
	.w2(32'h3bb47208),
	.w3(32'h39c5f652),
	.w4(32'h3bd1ea6a),
	.w5(32'h3c124747),
	.w6(32'h3bbd926b),
	.w7(32'h3ba662de),
	.w8(32'h3a9cc211),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b84298a),
	.w1(32'h3a6ba7bb),
	.w2(32'h3ae882ef),
	.w3(32'h3b961cef),
	.w4(32'h3a4b2f97),
	.w5(32'h3a2fbeb3),
	.w6(32'h3a506aeb),
	.w7(32'h3aa6dbcb),
	.w8(32'h3887f2af),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d14c9d),
	.w1(32'hb898d56e),
	.w2(32'h3946d222),
	.w3(32'hb992602a),
	.w4(32'hb904e053),
	.w5(32'hba105652),
	.w6(32'hb948de39),
	.w7(32'hb9828616),
	.w8(32'hba781744),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a67aae),
	.w1(32'hbb2d03ed),
	.w2(32'hba82b9ec),
	.w3(32'hba2bf120),
	.w4(32'hbb2c1e05),
	.w5(32'hbab626fc),
	.w6(32'hbb6b766c),
	.w7(32'hbb0a7d85),
	.w8(32'hba6d6591),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0e4779),
	.w1(32'hbb478da6),
	.w2(32'hbb8af32d),
	.w3(32'hba89f92b),
	.w4(32'hbb458eb7),
	.w5(32'hbb33716e),
	.w6(32'hbb57112f),
	.w7(32'hbb93cd17),
	.w8(32'hbaf81029),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb369e75),
	.w1(32'hba9583ba),
	.w2(32'hba0c5c61),
	.w3(32'hbabba34f),
	.w4(32'hba08c50d),
	.w5(32'hba1d5f27),
	.w6(32'hbac640da),
	.w7(32'hbaa0ed0a),
	.w8(32'hbb297e0c),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9d727a),
	.w1(32'hb553fdc4),
	.w2(32'h3a4c7ce4),
	.w3(32'hbb1944ca),
	.w4(32'h384b833f),
	.w5(32'hb8d73f83),
	.w6(32'hb8e044ae),
	.w7(32'h393ab1a8),
	.w8(32'hb9396501),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b44aaaf),
	.w1(32'hba66a66e),
	.w2(32'hbab6b5d3),
	.w3(32'h3ae4d3d6),
	.w4(32'hbb0e0b38),
	.w5(32'hbb0897c0),
	.w6(32'h3adb6f15),
	.w7(32'hba92da9f),
	.w8(32'hbaca6f23),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b154983),
	.w1(32'h3ac67cee),
	.w2(32'hba412b13),
	.w3(32'hba5e387b),
	.w4(32'hb9ae98c6),
	.w5(32'hbb6871c7),
	.w6(32'h3b0e7fc4),
	.w7(32'h3b1c0fc4),
	.w8(32'hbb3d0f10),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb09b718),
	.w1(32'h39a1c658),
	.w2(32'hbb031b8e),
	.w3(32'hbb372a75),
	.w4(32'h39fd83e2),
	.w5(32'hbb69a8a4),
	.w6(32'hba96c162),
	.w7(32'hb9033129),
	.w8(32'hbb2585d7),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3959f47a),
	.w1(32'h39c1bb83),
	.w2(32'h39de3db8),
	.w3(32'h3952cffa),
	.w4(32'h39936d29),
	.w5(32'h399de020),
	.w6(32'h3a4ddbcb),
	.w7(32'h39f5d818),
	.w8(32'hba31725f),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fc3a55),
	.w1(32'h3b0659ef),
	.w2(32'h3b1daec8),
	.w3(32'h39d626ba),
	.w4(32'h3b984d09),
	.w5(32'h3bd9e560),
	.w6(32'h3b91cf14),
	.w7(32'h3b764e6d),
	.w8(32'h3b6100a8),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b875d4d),
	.w1(32'h387f01dd),
	.w2(32'h395ce615),
	.w3(32'h3b9f4bc9),
	.w4(32'hba954077),
	.w5(32'hba88b5cc),
	.w6(32'hba48b874),
	.w7(32'hba1abdf5),
	.w8(32'hba85881c),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba67f080),
	.w1(32'h39b01330),
	.w2(32'h3919e379),
	.w3(32'hbaef9822),
	.w4(32'h39b269ac),
	.w5(32'hb9ad9601),
	.w6(32'hb9cd27e7),
	.w7(32'hb8278788),
	.w8(32'hbb0084f6),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8097ac),
	.w1(32'h3b47570d),
	.w2(32'h3b9e51a0),
	.w3(32'hbab59441),
	.w4(32'h3ad5ae0c),
	.w5(32'h3b5b5d3c),
	.w6(32'hba8e52d3),
	.w7(32'hbaa3ab6e),
	.w8(32'hb9b40d69),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b747428),
	.w1(32'h3ad97afe),
	.w2(32'h3a7c6984),
	.w3(32'h3ac3a1f1),
	.w4(32'h3aeefbb2),
	.w5(32'h3aa654ac),
	.w6(32'h3aafb956),
	.w7(32'hb8f081cb),
	.w8(32'hb78a11ed),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4273db),
	.w1(32'h38fb788b),
	.w2(32'hb972f753),
	.w3(32'h3a99f812),
	.w4(32'hbae1dcdf),
	.w5(32'hba23b318),
	.w6(32'hba36ba88),
	.w7(32'hbb3bc173),
	.w8(32'hbb1c3974),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac763a4),
	.w1(32'h3ad9afe6),
	.w2(32'h3a4f450e),
	.w3(32'hb9b8325b),
	.w4(32'hba5bf02a),
	.w5(32'h3a3c699e),
	.w6(32'h39e9cda9),
	.w7(32'h3a3374d2),
	.w8(32'h3a416789),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8adf9e6),
	.w1(32'h3b1861a5),
	.w2(32'h3baffa61),
	.w3(32'h39cd9992),
	.w4(32'h390ab440),
	.w5(32'h3b7e4756),
	.w6(32'h3ac71ddc),
	.w7(32'h3b4c2c10),
	.w8(32'hba00e2f0),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b31bfb8),
	.w1(32'hba8f7ffb),
	.w2(32'hb93fd0c6),
	.w3(32'hba9c23b2),
	.w4(32'hba1d74e2),
	.w5(32'hb9ca2a84),
	.w6(32'hbabd342b),
	.w7(32'hba675608),
	.w8(32'hbad355f2),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad2240d),
	.w1(32'h3a82676b),
	.w2(32'h3a06cf29),
	.w3(32'hbb1b6dd8),
	.w4(32'hb8c11249),
	.w5(32'hb9224fc8),
	.w6(32'hb93f6d8a),
	.w7(32'hba498e6a),
	.w8(32'h3a170fec),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f6ac3f),
	.w1(32'h39f09c8e),
	.w2(32'hb98bccfd),
	.w3(32'hb9507a45),
	.w4(32'hb9c028f8),
	.w5(32'hba1fe857),
	.w6(32'hb9cabf09),
	.w7(32'hba769784),
	.w8(32'hbadca088),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399e9217),
	.w1(32'h3b3368c5),
	.w2(32'h3a24c05e),
	.w3(32'hb9a276b0),
	.w4(32'h3b244425),
	.w5(32'h39da637b),
	.w6(32'h3b4e8ee8),
	.w7(32'h3a951049),
	.w8(32'h3a5aec9b),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a754324),
	.w1(32'h3a6e4103),
	.w2(32'h3b005aaf),
	.w3(32'h3a55b415),
	.w4(32'h3a3da246),
	.w5(32'h3a9f20af),
	.w6(32'h3a0138af),
	.w7(32'h3a34449b),
	.w8(32'h39e3038d),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b413f6a),
	.w1(32'h3ab29981),
	.w2(32'h3a990c51),
	.w3(32'hb9785bb3),
	.w4(32'hba957a64),
	.w5(32'h39c52b31),
	.w6(32'hb91c8590),
	.w7(32'hbaa3f0f2),
	.w8(32'h39693de2),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a58879f),
	.w1(32'hbaf065dc),
	.w2(32'h399c2436),
	.w3(32'h399fe252),
	.w4(32'hba0a4849),
	.w5(32'h3aede16c),
	.w6(32'hbb16e7a4),
	.w7(32'h39175d6f),
	.w8(32'hba820479),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7fe027),
	.w1(32'h397b15be),
	.w2(32'hb894f17f),
	.w3(32'h3927e7fa),
	.w4(32'h3ac44596),
	.w5(32'h3a9bc1b4),
	.w6(32'h3b777a84),
	.w7(32'h3b49515b),
	.w8(32'h3b644ad1),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5a2f89),
	.w1(32'hba38978a),
	.w2(32'hba724af1),
	.w3(32'h3aabe008),
	.w4(32'hb9ad4736),
	.w5(32'h36ae1c05),
	.w6(32'h3a030647),
	.w7(32'hb96f7c59),
	.w8(32'hba875c10),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacb2f56),
	.w1(32'h39df3180),
	.w2(32'hb914789a),
	.w3(32'hba4bb7f6),
	.w4(32'hb8974d5d),
	.w5(32'hb9f147ad),
	.w6(32'h3a69cfd1),
	.w7(32'hb99bf8eb),
	.w8(32'hba6c5f63),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba51ca71),
	.w1(32'h3aa9a7d3),
	.w2(32'h3a0e9f9a),
	.w3(32'hba16d276),
	.w4(32'h3aab9191),
	.w5(32'h39fec068),
	.w6(32'h3abc4d49),
	.w7(32'h3a40b004),
	.w8(32'hba1f5243),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398b18bc),
	.w1(32'hb991a393),
	.w2(32'hb9c2d4cc),
	.w3(32'h3a21722e),
	.w4(32'h385adc70),
	.w5(32'hba33d028),
	.w6(32'h395256c0),
	.w7(32'hb88bf5fd),
	.w8(32'hb8f29604),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37d2d8f5),
	.w1(32'h3aaa6c7f),
	.w2(32'h3b0b1a62),
	.w3(32'hba60db65),
	.w4(32'h3a2c1f15),
	.w5(32'h3ab4ad8b),
	.w6(32'hb9ca4d6f),
	.w7(32'hb8864dfe),
	.w8(32'h395505ad),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ace86c4),
	.w1(32'h39d1972f),
	.w2(32'h3a3b9e6d),
	.w3(32'h3a3c5ece),
	.w4(32'h3a7740ee),
	.w5(32'h3a268903),
	.w6(32'h39bf803c),
	.w7(32'h39ef9dea),
	.w8(32'h3a574679),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a322ce),
	.w1(32'hbacd5e78),
	.w2(32'hbb3d96f2),
	.w3(32'h39c34738),
	.w4(32'hb9b13393),
	.w5(32'hbab64f60),
	.w6(32'hbb302796),
	.w7(32'hbb49c1b5),
	.w8(32'h3a794b1b),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7782f6),
	.w1(32'h3a254395),
	.w2(32'h3a08914c),
	.w3(32'h398198eb),
	.w4(32'h3a56c0c5),
	.w5(32'h3a2378ee),
	.w6(32'h38b415cc),
	.w7(32'hb95a37ac),
	.w8(32'hba1b9b98),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b4c87c),
	.w1(32'hb9b4df01),
	.w2(32'h39f081fa),
	.w3(32'hb9af8eda),
	.w4(32'hba1d1561),
	.w5(32'hb9412c70),
	.w6(32'hb9de50f3),
	.w7(32'h39bceaa3),
	.w8(32'h39a868e0),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a00ab7c),
	.w1(32'h3a9e5322),
	.w2(32'h3a08125b),
	.w3(32'h39c5cf0b),
	.w4(32'hb926f3e8),
	.w5(32'hb9c1f6e7),
	.w6(32'h3a509c89),
	.w7(32'hb7cc93cc),
	.w8(32'hba8bad0b),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39867977),
	.w1(32'h3ac7c45a),
	.w2(32'h3b3417d7),
	.w3(32'hbaa86956),
	.w4(32'h3a28f39e),
	.w5(32'h3b2186bf),
	.w6(32'h39fe5d47),
	.w7(32'h393f2555),
	.w8(32'h3b1b9773),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b35e519),
	.w1(32'h3bf185be),
	.w2(32'h3c160edc),
	.w3(32'h3b1a0608),
	.w4(32'h3bd1fa96),
	.w5(32'h3c27fcc0),
	.w6(32'h3bd64025),
	.w7(32'h3bd92723),
	.w8(32'h3b71805e),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c07e224),
	.w1(32'h38949b66),
	.w2(32'h3a3dcb16),
	.w3(32'h3bbc2630),
	.w4(32'hba921ffc),
	.w5(32'hba81edeb),
	.w6(32'hbaa9856a),
	.w7(32'hba4d9f63),
	.w8(32'hba87f11b),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7036c8),
	.w1(32'h3abbdde3),
	.w2(32'hba75dbde),
	.w3(32'h38b9112b),
	.w4(32'hb98c07bb),
	.w5(32'hbb10b795),
	.w6(32'h3a63bce7),
	.w7(32'hba9afc3c),
	.w8(32'hbb8ee0b0),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba66a558),
	.w1(32'h39cf31f1),
	.w2(32'h3a1e7f1b),
	.w3(32'hba11c72b),
	.w4(32'hb8984748),
	.w5(32'h390a43d9),
	.w6(32'h380b9286),
	.w7(32'h38496694),
	.w8(32'hba8a4a21),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e5fd44),
	.w1(32'hb8e83b4b),
	.w2(32'hb99b5521),
	.w3(32'hba7f996f),
	.w4(32'hba1639be),
	.w5(32'hba8a1b1f),
	.w6(32'h3974cc3c),
	.w7(32'hb921995a),
	.w8(32'hb9b405da),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba26638b),
	.w1(32'h38b9fa9e),
	.w2(32'h3871a5dc),
	.w3(32'hba6a5a17),
	.w4(32'hb8ab27b3),
	.w5(32'hba048fae),
	.w6(32'h39a523f7),
	.w7(32'hb9196de1),
	.w8(32'h3712c83a),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99d4a1f),
	.w1(32'h38267970),
	.w2(32'h3a9a06ac),
	.w3(32'hba6eff8f),
	.w4(32'hba5aac65),
	.w5(32'hb9dcb99d),
	.w6(32'hba5027b5),
	.w7(32'hb9aa9f91),
	.w8(32'hba5e54b2),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96879cd),
	.w1(32'h3af7165b),
	.w2(32'h3aaf54c5),
	.w3(32'hbae1fedc),
	.w4(32'h3aa7a3c5),
	.w5(32'h3a044bb8),
	.w6(32'h3ac6594b),
	.w7(32'h3a79fbdb),
	.w8(32'h3a4bf02f),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab48dcb),
	.w1(32'h39ef0ffb),
	.w2(32'hb714cf4a),
	.w3(32'hb870aadc),
	.w4(32'hbaa1fe88),
	.w5(32'hb9f00c2f),
	.w6(32'hb9ca209c),
	.w7(32'h37f88e74),
	.w8(32'hb958a08f),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba676397),
	.w1(32'h3a09267a),
	.w2(32'h3b0f6b9d),
	.w3(32'hbabb1ccc),
	.w4(32'hba089a33),
	.w5(32'hb9ff991c),
	.w6(32'hba5a4748),
	.w7(32'hb9d9ca50),
	.w8(32'h3a1373e9),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5daf7c),
	.w1(32'h39b92076),
	.w2(32'h3918f62e),
	.w3(32'hb8d6bde1),
	.w4(32'h394f2f94),
	.w5(32'h3a354dc8),
	.w6(32'h387195e8),
	.w7(32'hba0b4563),
	.w8(32'hba4e65bc),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a90c31b),
	.w1(32'hbb172ea6),
	.w2(32'h3b00bc2b),
	.w3(32'h390c9b5c),
	.w4(32'hb9dfad61),
	.w5(32'h3b74ec5d),
	.w6(32'hbb8354c4),
	.w7(32'h39c70bf7),
	.w8(32'hbb1dc3ab),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7b653b),
	.w1(32'h3ab50703),
	.w2(32'h3b235143),
	.w3(32'h39d2e1dc),
	.w4(32'h3a33eff3),
	.w5(32'h39c8296b),
	.w6(32'h3a2de0f3),
	.w7(32'h3a6e947c),
	.w8(32'hb8bb1ae4),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a55b6f9),
	.w1(32'h3ba1e9b9),
	.w2(32'h3b57d990),
	.w3(32'h392d6938),
	.w4(32'h3b4223e9),
	.w5(32'h3b4208fa),
	.w6(32'h3c05ff85),
	.w7(32'h3b9b8904),
	.w8(32'h3bdd26a2),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd274ad),
	.w1(32'h3a63aa81),
	.w2(32'h3a721b30),
	.w3(32'h3b58e048),
	.w4(32'hb8f72d4c),
	.w5(32'h3930d28b),
	.w6(32'h39621cb8),
	.w7(32'hb9eeca8d),
	.w8(32'hb9ce73a2),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb842d4e0),
	.w1(32'h3989c93a),
	.w2(32'h3a445ad7),
	.w3(32'hba8184a0),
	.w4(32'hb9b6bcfe),
	.w5(32'hb882cad4),
	.w6(32'h39831db1),
	.w7(32'h3a1b210e),
	.w8(32'hb70da129),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393acdc7),
	.w1(32'h3a959e2e),
	.w2(32'h3a5d99e2),
	.w3(32'hba477945),
	.w4(32'h3aa18b35),
	.w5(32'h3a2be608),
	.w6(32'h3a6571eb),
	.w7(32'h39de1c33),
	.w8(32'hb5901d2b),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39994338),
	.w1(32'h3b25e858),
	.w2(32'h3b675a3c),
	.w3(32'h38e165bf),
	.w4(32'hbb4912af),
	.w5(32'hba65e7e5),
	.w6(32'h3a4fdee3),
	.w7(32'h3b025d27),
	.w8(32'hb9f44237),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7cba9e),
	.w1(32'hba2e8421),
	.w2(32'hba08e02c),
	.w3(32'hbb6733ab),
	.w4(32'hba394e36),
	.w5(32'hb9116b54),
	.w6(32'h384ce351),
	.w7(32'h38d46e71),
	.w8(32'hba070d95),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb950aa36),
	.w1(32'h38a5463b),
	.w2(32'hba9406bf),
	.w3(32'hba2e3bee),
	.w4(32'hba197236),
	.w5(32'hba9edbf0),
	.w6(32'hb9f2f722),
	.w7(32'hba87ca36),
	.w8(32'hbb2b3868),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac69f28),
	.w1(32'h3a67cc8f),
	.w2(32'h3aa956de),
	.w3(32'hba8b6e72),
	.w4(32'h3a4bab1f),
	.w5(32'h3986b1ee),
	.w6(32'h3a995deb),
	.w7(32'h3aaefab0),
	.w8(32'hb8bc8d9a),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a56a31d),
	.w1(32'hbac9d1e2),
	.w2(32'hba5ed11b),
	.w3(32'hb99347a8),
	.w4(32'hba4be257),
	.w5(32'h3a6f2a43),
	.w6(32'hbaab5556),
	.w7(32'hbabc4be2),
	.w8(32'hbaf00729),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2693c4),
	.w1(32'h3acdf74f),
	.w2(32'h3b3d7238),
	.w3(32'hbaa7dfc5),
	.w4(32'h39c1a90c),
	.w5(32'h3a4f6469),
	.w6(32'h390da70f),
	.w7(32'h3a389b3d),
	.w8(32'hb94adbb9),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96ba1a2),
	.w1(32'h3ae966b5),
	.w2(32'h3acf844f),
	.w3(32'hba42cf22),
	.w4(32'h3a1d976c),
	.w5(32'hba885c86),
	.w6(32'h3a988cdc),
	.w7(32'h3ad0b882),
	.w8(32'hba99c44c),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b34a441),
	.w1(32'hb8b46072),
	.w2(32'h3a50af14),
	.w3(32'hba6f46ab),
	.w4(32'hbb0a77fb),
	.w5(32'hb7964e8a),
	.w6(32'hbaefdca6),
	.w7(32'hbb359397),
	.w8(32'hbb1fdc88),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b4fb51),
	.w1(32'h3900fc6d),
	.w2(32'h39e26002),
	.w3(32'hb9be2938),
	.w4(32'hb88c2ace),
	.w5(32'hba207c71),
	.w6(32'h3a825dbe),
	.w7(32'h3a889510),
	.w8(32'hba37cb29),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b27afe8),
	.w1(32'h3bcc7091),
	.w2(32'h3b6e66c7),
	.w3(32'hbae700d1),
	.w4(32'h3b20d294),
	.w5(32'h39a1bbee),
	.w6(32'h3bb030f4),
	.w7(32'h3b3e8cd5),
	.w8(32'h3ba91296),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc22cb2),
	.w1(32'h37201f69),
	.w2(32'hb93f4a0b),
	.w3(32'h3b34dc25),
	.w4(32'hba7aae9f),
	.w5(32'hb9c4d547),
	.w6(32'hba881e33),
	.w7(32'hbaa129d8),
	.w8(32'hbb0e852c),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39de0859),
	.w1(32'h3b03a642),
	.w2(32'h3a9ab449),
	.w3(32'hb787b556),
	.w4(32'h3a95229d),
	.w5(32'hb9cffafd),
	.w6(32'h3b4d52ee),
	.w7(32'h3b19648e),
	.w8(32'h38612d52),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac33915),
	.w1(32'h3b60c8cb),
	.w2(32'h3bc75427),
	.w3(32'h3a96e78b),
	.w4(32'h3ac431e9),
	.w5(32'h3bd56ea6),
	.w6(32'h3a1df65a),
	.w7(32'h3b736738),
	.w8(32'h3b0c2059),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be1ab19),
	.w1(32'hba2ca0fe),
	.w2(32'h39af76dd),
	.w3(32'h3b559023),
	.w4(32'hbae3cf74),
	.w5(32'hb8829854),
	.w6(32'hbb551a8c),
	.w7(32'hbb9491cd),
	.w8(32'hbb2c0a4c),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9674fe),
	.w1(32'h3a0b7504),
	.w2(32'h3aa0828c),
	.w3(32'hbb48d26a),
	.w4(32'hbaa7ebd5),
	.w5(32'hba3b3c2f),
	.w6(32'hbb2f56c6),
	.w7(32'hba083890),
	.w8(32'hba998563),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c39a4b),
	.w1(32'h39aedaf0),
	.w2(32'h3b1abd32),
	.w3(32'hba3d8cc9),
	.w4(32'hb8f29d8e),
	.w5(32'h3adef5df),
	.w6(32'h3ad7ccbc),
	.w7(32'h3988d99d),
	.w8(32'h38b7dc6e),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3becaa1c),
	.w1(32'h3ac39d4d),
	.w2(32'hbb8b2cf7),
	.w3(32'h3bcb63e5),
	.w4(32'hbb2b1ee0),
	.w5(32'hbbc90759),
	.w6(32'h39759241),
	.w7(32'hbb93e0fa),
	.w8(32'hbc0c8e5d),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1459ee),
	.w1(32'h385c171b),
	.w2(32'hbae50200),
	.w3(32'hba123f80),
	.w4(32'hbb06c96d),
	.w5(32'hbb0a2897),
	.w6(32'h3a49b9d8),
	.w7(32'hba9473da),
	.w8(32'h3a56995f),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b059b62),
	.w1(32'h3a8acac0),
	.w2(32'h3a708eb7),
	.w3(32'h3af03202),
	.w4(32'hba5736b4),
	.w5(32'hba958d06),
	.w6(32'h3a289f0d),
	.w7(32'hba557962),
	.w8(32'hb91babe0),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ffe967),
	.w1(32'h3a3acce5),
	.w2(32'h39757680),
	.w3(32'hba633ca4),
	.w4(32'h39ffec68),
	.w5(32'hb999dcf4),
	.w6(32'hba191724),
	.w7(32'hb9d3589a),
	.w8(32'h3733d695),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaf066c),
	.w1(32'h3a461ae1),
	.w2(32'h39e22d37),
	.w3(32'hb916d236),
	.w4(32'hba98fb9a),
	.w5(32'hbadcec4e),
	.w6(32'h3a52d098),
	.w7(32'hb9e66570),
	.w8(32'h3943cc01),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e7d1a2),
	.w1(32'hbaaca935),
	.w2(32'hb9245ba8),
	.w3(32'hba2f3db1),
	.w4(32'hb9b4dab1),
	.w5(32'h39b421c0),
	.w6(32'hba15a830),
	.w7(32'hb8a9434f),
	.w8(32'h3960476b),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9b24c3),
	.w1(32'h3a24641b),
	.w2(32'h3a1a5121),
	.w3(32'hba9165dc),
	.w4(32'hb7c45ec9),
	.w5(32'hb8f00ead),
	.w6(32'hb920c2ef),
	.w7(32'h38b28ef4),
	.w8(32'hba0513c3),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f3d5c6),
	.w1(32'h3b35c8e2),
	.w2(32'h3b8d333f),
	.w3(32'hba7ee373),
	.w4(32'h3a9cde52),
	.w5(32'h3a9c599b),
	.w6(32'h3ac9d388),
	.w7(32'h3b1a2b9b),
	.w8(32'hb9847760),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b44b7b6),
	.w1(32'hb9bf6d6f),
	.w2(32'h3a3a5b4f),
	.w3(32'hba8cd930),
	.w4(32'hbaa4a7c4),
	.w5(32'hb89c8777),
	.w6(32'hbaa2391c),
	.w7(32'hbb1c86ad),
	.w8(32'hb91191fc),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3add15bb),
	.w1(32'h3950cb15),
	.w2(32'hb9562dee),
	.w3(32'hb8b95f05),
	.w4(32'hbabe7253),
	.w5(32'hba6a15e0),
	.w6(32'hba774daa),
	.w7(32'hbb1751f5),
	.w8(32'hbb1dc27d),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39882f47),
	.w1(32'h3a729e73),
	.w2(32'hba272d84),
	.w3(32'h38322321),
	.w4(32'h39e85078),
	.w5(32'hbb024833),
	.w6(32'h39cdad13),
	.w7(32'hb9dac0da),
	.w8(32'hbacb6de2),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8e1ce2),
	.w1(32'h3ab34710),
	.w2(32'hb97103dc),
	.w3(32'hb91abc57),
	.w4(32'h3b441f98),
	.w5(32'h38efcb1f),
	.w6(32'hba6fa1b0),
	.w7(32'hbab48da9),
	.w8(32'h3a242f3d),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99c1fc6),
	.w1(32'hba511bc1),
	.w2(32'hba8bece3),
	.w3(32'hbad4ac8f),
	.w4(32'hba82bc5c),
	.w5(32'hbb114a83),
	.w6(32'hb9718540),
	.w7(32'hba59dd91),
	.w8(32'hbaa68ff0),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0f39ff),
	.w1(32'hb936c4d1),
	.w2(32'h3a021e07),
	.w3(32'h38d187ea),
	.w4(32'h38f627ef),
	.w5(32'h39921d53),
	.w6(32'h38f81747),
	.w7(32'hba1b4a7e),
	.w8(32'hbaa07e21),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8dcead),
	.w1(32'hbb03b2b0),
	.w2(32'hbb0f6df7),
	.w3(32'h399f6166),
	.w4(32'hbae5bb3d),
	.w5(32'hbafd8759),
	.w6(32'hbac31b1e),
	.w7(32'hbb0f16ab),
	.w8(32'hba94dcb1),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaf0602),
	.w1(32'h3862d3cd),
	.w2(32'h3987308c),
	.w3(32'hbab086ac),
	.w4(32'h383f113f),
	.w5(32'hba57c618),
	.w6(32'h3997ba71),
	.w7(32'h3893594f),
	.w8(32'h3962104f),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h373d1de1),
	.w1(32'hb8da5f5b),
	.w2(32'h39b2042d),
	.w3(32'hba476ec3),
	.w4(32'hba0a8b67),
	.w5(32'hba47a411),
	.w6(32'h37413e40),
	.w7(32'hb8e70717),
	.w8(32'hb9044f11),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9501998),
	.w1(32'hb9a2613a),
	.w2(32'h392a82b5),
	.w3(32'hba36987b),
	.w4(32'hba0ad948),
	.w5(32'hba856839),
	.w6(32'hb8a97607),
	.w7(32'hb9227e06),
	.w8(32'hb903dc40),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba06ba48),
	.w1(32'h37e0dc0d),
	.w2(32'h39723c6a),
	.w3(32'hba86c1cf),
	.w4(32'h3a158fb6),
	.w5(32'h3a1702b8),
	.w6(32'h375be034),
	.w7(32'h3a8a1b2b),
	.w8(32'h39ef6601),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6947e1),
	.w1(32'hb98c9c48),
	.w2(32'h39609f92),
	.w3(32'h3798649b),
	.w4(32'hbac64c11),
	.w5(32'h393d5cef),
	.w6(32'h39cec7d3),
	.w7(32'hb9dbe047),
	.w8(32'hbacf5d01),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba39a0b1),
	.w1(32'hba2b7791),
	.w2(32'hb9aa5636),
	.w3(32'hb8853862),
	.w4(32'hba087723),
	.w5(32'hbaca5f57),
	.w6(32'hb68985dc),
	.w7(32'hb9dec260),
	.w8(32'hb98f599d),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395167d0),
	.w1(32'h39bb2084),
	.w2(32'h3a20aa6f),
	.w3(32'hbac1d624),
	.w4(32'h387dd69f),
	.w5(32'hb9206fbb),
	.w6(32'h3947d6de),
	.w7(32'hb99734ce),
	.w8(32'hba7dc69a),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1d26be),
	.w1(32'h3988e698),
	.w2(32'hba8082af),
	.w3(32'hba649515),
	.w4(32'h385d5e84),
	.w5(32'hbb054870),
	.w6(32'h3a7c2342),
	.w7(32'h39ca963a),
	.w8(32'hba540221),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3921ba64),
	.w1(32'hbaaf56a4),
	.w2(32'hbadeab0b),
	.w3(32'hb92557c9),
	.w4(32'hb9dcbbd4),
	.w5(32'hb9eadfde),
	.w6(32'hb8ff8445),
	.w7(32'h3a76550b),
	.w8(32'h39aa5c7c),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb02c7a5),
	.w1(32'h3a651866),
	.w2(32'h3aa0155b),
	.w3(32'hb997ec95),
	.w4(32'h39cb7b5e),
	.w5(32'hb8e3e6e3),
	.w6(32'h3a519fcf),
	.w7(32'h3a0872d6),
	.w8(32'h39815ecd),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa5eeb2),
	.w1(32'h3a986ee5),
	.w2(32'h3b014b4c),
	.w3(32'hb8a734b4),
	.w4(32'h3a328f78),
	.w5(32'hb8937961),
	.w6(32'h3a86c9ec),
	.w7(32'h3a6e9e53),
	.w8(32'hb8f4afdd),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a253178),
	.w1(32'hb960775b),
	.w2(32'hb8fbd0c1),
	.w3(32'hba70c58b),
	.w4(32'hb9f4e8ba),
	.w5(32'hb9a7c9b6),
	.w6(32'hb9beea22),
	.w7(32'hba2ae8bf),
	.w8(32'hb9e47cd7),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39842315),
	.w1(32'hb9dde201),
	.w2(32'h38adf059),
	.w3(32'hba801a1a),
	.w4(32'hba14c6b8),
	.w5(32'h3a2207ab),
	.w6(32'hb9904f81),
	.w7(32'hba370b1f),
	.w8(32'hb69cd387),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ae4359),
	.w1(32'hb8b01a4c),
	.w2(32'h3ad46bb5),
	.w3(32'hba555fb9),
	.w4(32'hbab3dc2c),
	.w5(32'h3a4a1a00),
	.w6(32'hba32b688),
	.w7(32'hbac21839),
	.w8(32'h37c519e5),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38573fa9),
	.w1(32'h38b64c16),
	.w2(32'h39081b43),
	.w3(32'hb8fe94a0),
	.w4(32'hb8a02d73),
	.w5(32'hb716661c),
	.w6(32'hb875d4bb),
	.w7(32'hb89a5006),
	.w8(32'hb82316d0),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b4efbe),
	.w1(32'hb764f604),
	.w2(32'hb38b04a0),
	.w3(32'hb88f679e),
	.w4(32'hb998ae78),
	.w5(32'hb9c75e53),
	.w6(32'hb93db7fd),
	.w7(32'hba060c6b),
	.w8(32'hb9d59461),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39498d44),
	.w1(32'h38ed29c0),
	.w2(32'hb881bdb5),
	.w3(32'h389ac8a5),
	.w4(32'h38a9373d),
	.w5(32'hb9324c3d),
	.w6(32'h3829d74c),
	.w7(32'h383f6f37),
	.w8(32'hb91a5164),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1fee55),
	.w1(32'h3801f5be),
	.w2(32'h391dbc3c),
	.w3(32'hb6fd0c48),
	.w4(32'hba07e2dd),
	.w5(32'hb867f30e),
	.w6(32'hba1af33b),
	.w7(32'hba752368),
	.w8(32'hb94f5e5e),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f94e7a),
	.w1(32'h3a1fa022),
	.w2(32'h3a51ea99),
	.w3(32'hba0cf587),
	.w4(32'hba10e1b1),
	.w5(32'h38862f8c),
	.w6(32'hbacec8ae),
	.w7(32'hba942aab),
	.w8(32'hb9572e7a),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a992287),
	.w1(32'h39a07f18),
	.w2(32'h3a852f53),
	.w3(32'hba0bbaea),
	.w4(32'hba3caede),
	.w5(32'h399a5707),
	.w6(32'hb99c37ec),
	.w7(32'hba25cf87),
	.w8(32'hb896cada),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2afaaf),
	.w1(32'h38b3f693),
	.w2(32'hba1d7216),
	.w3(32'h3a031c57),
	.w4(32'hb9655c7e),
	.w5(32'hba263e43),
	.w6(32'h38c36f85),
	.w7(32'hba4a0fca),
	.w8(32'hba68f348),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a69cb09),
	.w1(32'hb91108e1),
	.w2(32'hb6d5b838),
	.w3(32'h392ce3f5),
	.w4(32'hba369ba6),
	.w5(32'hba4302a4),
	.w6(32'hb5f63100),
	.w7(32'hba7543c1),
	.w8(32'hba07486a),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a60e0e1),
	.w1(32'h39f4df3f),
	.w2(32'h3a2823a1),
	.w3(32'hb907471d),
	.w4(32'hba07e785),
	.w5(32'hb8bfba5c),
	.w6(32'hb907512b),
	.w7(32'hba37d480),
	.w8(32'hb9c0d2c9),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e21ece),
	.w1(32'hb99d6040),
	.w2(32'hba2deb10),
	.w3(32'hb92986ee),
	.w4(32'hba396172),
	.w5(32'hba5e950e),
	.w6(32'h38c4b209),
	.w7(32'hb9eb402a),
	.w8(32'hba4efbb2),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae2636a),
	.w1(32'h39b8ddad),
	.w2(32'h3a144d05),
	.w3(32'h3a3cceca),
	.w4(32'hb9e7ca51),
	.w5(32'h39547911),
	.w6(32'h38b87dcb),
	.w7(32'hba8f9aaf),
	.w8(32'hb946d310),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bb9a0c),
	.w1(32'h38c45426),
	.w2(32'h390a1c1b),
	.w3(32'h3933edc9),
	.w4(32'hb942c309),
	.w5(32'h38c1d001),
	.w6(32'hb8a48b1f),
	.w7(32'hb9e7edac),
	.w8(32'hb8e5a9c1),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac28482),
	.w1(32'h3a2cc2aa),
	.w2(32'hbacb5d0d),
	.w3(32'h396deb91),
	.w4(32'hb699de00),
	.w5(32'hbae79673),
	.w6(32'h3a3526a2),
	.w7(32'h3a30a6fe),
	.w8(32'hba9dbc1e),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d0c147),
	.w1(32'hb831b190),
	.w2(32'h385d1650),
	.w3(32'h3925d12b),
	.w4(32'hb9d34e7c),
	.w5(32'hb9971b53),
	.w6(32'hb994d1c1),
	.w7(32'hb9f7e3fe),
	.w8(32'h38543187),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb79437c4),
	.w1(32'h36806fbb),
	.w2(32'h378eaab1),
	.w3(32'hb5c254a1),
	.w4(32'h36c04f54),
	.w5(32'h37c3977f),
	.w6(32'h37463e1d),
	.w7(32'hb780901d),
	.w8(32'h37baa728),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7c25b34),
	.w1(32'h351ebdd6),
	.w2(32'hb83565b5),
	.w3(32'hb72c51ab),
	.w4(32'hb7416c45),
	.w5(32'hb82d2822),
	.w6(32'h380501b5),
	.w7(32'h37caf793),
	.w8(32'hb81900ff),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389dd1d3),
	.w1(32'h3910b5a7),
	.w2(32'h376fabfa),
	.w3(32'h3668d088),
	.w4(32'hb91f8388),
	.w5(32'hb8ddc546),
	.w6(32'h3917c57d),
	.w7(32'h38fcbc50),
	.w8(32'hb8100c6c),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9a7300),
	.w1(32'h391f1bfb),
	.w2(32'hba59b007),
	.w3(32'h3a2ec628),
	.w4(32'hb8865a87),
	.w5(32'hba864198),
	.w6(32'h3a149d72),
	.w7(32'h39bfffd3),
	.w8(32'hb9d31ab6),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0306d7),
	.w1(32'h3a56a14d),
	.w2(32'h3aa6daa6),
	.w3(32'hb9cfe5bb),
	.w4(32'hb9b5ecfb),
	.w5(32'h3a0d81b6),
	.w6(32'hbaa3f21c),
	.w7(32'hba3031b8),
	.w8(32'h38d6e5c4),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7a09a71),
	.w1(32'h384768f1),
	.w2(32'hb7b51433),
	.w3(32'hb818432a),
	.w4(32'h37e99f0a),
	.w5(32'hb6f80908),
	.w6(32'hb5da0f86),
	.w7(32'hb72663eb),
	.w8(32'h37ed4823),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab6caae),
	.w1(32'h3a26eadc),
	.w2(32'h3aa6df62),
	.w3(32'hb883594a),
	.w4(32'hba5e5c4f),
	.w5(32'h3a1feedf),
	.w6(32'hba8b8b8d),
	.w7(32'hbac02905),
	.w8(32'h3778b2e1),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba421bcc),
	.w1(32'hba880a3a),
	.w2(32'hb84ce185),
	.w3(32'hbab8c155),
	.w4(32'hbacb31ed),
	.w5(32'h3a05034b),
	.w6(32'hba946443),
	.w7(32'hbac2fee4),
	.w8(32'h3a59a31b),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa3d3bf),
	.w1(32'hb9239128),
	.w2(32'hb81c8b8b),
	.w3(32'h3a76f596),
	.w4(32'hba2cef43),
	.w5(32'hb9f67928),
	.w6(32'h39b2d750),
	.w7(32'hba829e9f),
	.w8(32'hba4aa036),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a008a3f),
	.w1(32'h3a9d9e18),
	.w2(32'h3a0a5147),
	.w3(32'hba1390ac),
	.w4(32'hb82ec6e7),
	.w5(32'hba0eab9f),
	.w6(32'h39bd2782),
	.w7(32'h39aab116),
	.w8(32'hb93e3236),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398cb893),
	.w1(32'h39ac1fa4),
	.w2(32'hb96e6e7c),
	.w3(32'hb9db210a),
	.w4(32'hb9c96552),
	.w5(32'hb986f8fc),
	.w6(32'hb9b6e637),
	.w7(32'h3657cbfd),
	.w8(32'hb809a650),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a200acb),
	.w1(32'h3a272d13),
	.w2(32'hba090222),
	.w3(32'h390d07f0),
	.w4(32'h38d98b0b),
	.w5(32'hb997899a),
	.w6(32'hba0a2f8b),
	.w7(32'hba4e0f0e),
	.w8(32'hb9ffdcf4),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b074f92),
	.w1(32'h39424c6a),
	.w2(32'hb8461d81),
	.w3(32'h3a779a0c),
	.w4(32'hb9d23962),
	.w5(32'hb987aded),
	.w6(32'h394d763a),
	.w7(32'hbaa2d509),
	.w8(32'hba30347b),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0b58fb),
	.w1(32'h3a6da372),
	.w2(32'h39f69d14),
	.w3(32'hba8c7608),
	.w4(32'hb896fa60),
	.w5(32'hb987b7fc),
	.w6(32'hba809221),
	.w7(32'h39dccf6c),
	.w8(32'h38e75d16),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d76405),
	.w1(32'hb920ee58),
	.w2(32'hba572656),
	.w3(32'hb9bd0f28),
	.w4(32'hb57045e8),
	.w5(32'hba526425),
	.w6(32'hb943aa38),
	.w7(32'h38eab057),
	.w8(32'hba3055c6),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393d1fea),
	.w1(32'h397f5933),
	.w2(32'h399e33b0),
	.w3(32'hb813f09d),
	.w4(32'h38bb16c1),
	.w5(32'h39002d9e),
	.w6(32'h3877e71c),
	.w7(32'hb6d135d9),
	.w8(32'h38142ffd),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h381cb4d8),
	.w1(32'h38146581),
	.w2(32'h376b9410),
	.w3(32'h378f6808),
	.w4(32'h38325e51),
	.w5(32'h37abe8ef),
	.w6(32'h3685fa7b),
	.w7(32'h3803b698),
	.w8(32'h3787a619),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a89f4bd),
	.w1(32'h39f1acc3),
	.w2(32'h39d0e72a),
	.w3(32'h391f3438),
	.w4(32'hb9c07395),
	.w5(32'hb9cd4606),
	.w6(32'hb9ab0d65),
	.w7(32'hba875e49),
	.w8(32'hba3ce7ac),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3944f259),
	.w1(32'h3984d3ab),
	.w2(32'h39257b84),
	.w3(32'h3892c21b),
	.w4(32'h39042b83),
	.w5(32'h389e9a80),
	.w6(32'h396b5514),
	.w7(32'h38a45d25),
	.w8(32'hb88facf8),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1c7432),
	.w1(32'hb84b09d2),
	.w2(32'h397f3913),
	.w3(32'h395ea892),
	.w4(32'hb9c6cb57),
	.w5(32'h38148b0e),
	.w6(32'h39e2fa19),
	.w7(32'hba2767d6),
	.w8(32'hb9be9ec0),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399caf21),
	.w1(32'hb91750cb),
	.w2(32'hb97d2af5),
	.w3(32'h39a48ec6),
	.w4(32'h395720a5),
	.w5(32'hb95259cf),
	.w6(32'h3994a55d),
	.w7(32'h39ef2910),
	.w8(32'hb98e83bf),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab7ead6),
	.w1(32'h3875c3a5),
	.w2(32'hb88533de),
	.w3(32'hbb10d057),
	.w4(32'hb804273c),
	.w5(32'h3846d78b),
	.w6(32'hbaec25e0),
	.w7(32'hb9f32c78),
	.w8(32'hb6d0e94a),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb912a0b7),
	.w1(32'h3880cfa3),
	.w2(32'h391e6f41),
	.w3(32'hb8a0583f),
	.w4(32'h383263c5),
	.w5(32'h38eda031),
	.w6(32'hb943a93c),
	.w7(32'hb7a80858),
	.w8(32'h38475760),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9539912),
	.w1(32'hb7a4f379),
	.w2(32'hb79e1220),
	.w3(32'hb9aed047),
	.w4(32'hb90b1209),
	.w5(32'hb8c411c3),
	.w6(32'hb9dd5333),
	.w7(32'hb9188ae7),
	.w8(32'hb895e2d4),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa1df03),
	.w1(32'h3a041be4),
	.w2(32'hb926c0dc),
	.w3(32'h39f96ee6),
	.w4(32'hba5c587b),
	.w5(32'hbac0acff),
	.w6(32'h39fe2ffe),
	.w7(32'hbaa6050a),
	.w8(32'hbb17e3c2),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0248fc),
	.w1(32'hb9134049),
	.w2(32'h38d4733a),
	.w3(32'h3a7ef91f),
	.w4(32'hba987a3b),
	.w5(32'h394f79e2),
	.w6(32'h3a2caa99),
	.w7(32'hbac7fec2),
	.w8(32'hb8288ca7),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4c2adb),
	.w1(32'hb9639f40),
	.w2(32'hba040e56),
	.w3(32'hba48f33f),
	.w4(32'hb8bf839d),
	.w5(32'hb9b4184d),
	.w6(32'hb9e7078a),
	.w7(32'h39101d9a),
	.w8(32'hb9e03ffd),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a975117),
	.w1(32'hba4f3e2f),
	.w2(32'hbaa96c30),
	.w3(32'h3ab53d3f),
	.w4(32'hb9e7bdf3),
	.w5(32'hb9ab824f),
	.w6(32'hb95c86a4),
	.w7(32'hbaeb37e7),
	.w8(32'hba77210a),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d6293b),
	.w1(32'h3892b3b2),
	.w2(32'h39990cdd),
	.w3(32'hb92c426a),
	.w4(32'hb91e979f),
	.w5(32'h395e6e31),
	.w6(32'hb9d71d35),
	.w7(32'hb91f3993),
	.w8(32'h377e75bc),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4060f0),
	.w1(32'h3a36f96b),
	.w2(32'h3a64056f),
	.w3(32'hb926a6b0),
	.w4(32'hb99fc73d),
	.w5(32'h3942847d),
	.w6(32'hba1c5715),
	.w7(32'hba543079),
	.w8(32'hb9429727),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa464c6),
	.w1(32'h3ab4f380),
	.w2(32'h3a881461),
	.w3(32'h3938a812),
	.w4(32'h388c479a),
	.w5(32'hb958a2e4),
	.w6(32'hba233984),
	.w7(32'hba1531ef),
	.w8(32'hb9f8b891),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2cb80e),
	.w1(32'h3a2bcd52),
	.w2(32'h3a89cc53),
	.w3(32'h3a6d9be1),
	.w4(32'hba5ce9d4),
	.w5(32'h39a6ad2a),
	.w6(32'hba498db2),
	.w7(32'hbb1ea58f),
	.w8(32'hb9a0e227),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388f3be0),
	.w1(32'h39893fff),
	.w2(32'h399e3a3f),
	.w3(32'h39affea4),
	.w4(32'h396ec83d),
	.w5(32'h386ad3d7),
	.w6(32'h3a18b7c9),
	.w7(32'h39b2bb6b),
	.w8(32'hb9c144c5),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1cac2c),
	.w1(32'h38505b65),
	.w2(32'h396d9340),
	.w3(32'h3966891f),
	.w4(32'hba0018a9),
	.w5(32'h36a128b4),
	.w6(32'hb82b311e),
	.w7(32'hb9c882d7),
	.w8(32'hb84c1954),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7587518),
	.w1(32'hb74d0cb9),
	.w2(32'hb7c17176),
	.w3(32'hb7cb200a),
	.w4(32'h36304254),
	.w5(32'hb6f35041),
	.w6(32'hb80e8aee),
	.w7(32'hb779fbc8),
	.w8(32'h37336d69),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397c54d6),
	.w1(32'h38925b70),
	.w2(32'hb908552c),
	.w3(32'hb8cc17f9),
	.w4(32'hb90e91cf),
	.w5(32'hb98c0d6e),
	.w6(32'hb9757557),
	.w7(32'hb995289b),
	.w8(32'hb9bf33cb),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ba9a21),
	.w1(32'hb75a4c15),
	.w2(32'hb98cab32),
	.w3(32'h39190dd5),
	.w4(32'h386767f7),
	.w5(32'hb9986f7f),
	.w6(32'h38a43cd8),
	.w7(32'h37f9db64),
	.w8(32'hb985477a),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a16604e),
	.w1(32'h39564b86),
	.w2(32'h396d99ab),
	.w3(32'hb945f419),
	.w4(32'hb9cb94ec),
	.w5(32'hb905a4ed),
	.w6(32'hba25fbf4),
	.w7(32'hba2b31d2),
	.w8(32'hb98c5c26),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7101382),
	.w1(32'h36d6ef27),
	.w2(32'hb749a10c),
	.w3(32'hb5eab744),
	.w4(32'h37172454),
	.w5(32'hb5eda5a4),
	.w6(32'h3703ca9e),
	.w7(32'h3682aa3b),
	.w8(32'h37de9570),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39109a89),
	.w1(32'h38df438b),
	.w2(32'h388b77db),
	.w3(32'hb7403648),
	.w4(32'hb8218e01),
	.w5(32'hb8cec40a),
	.w6(32'hb87b5f75),
	.w7(32'hb8cf9791),
	.w8(32'hb919ca98),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7c15343),
	.w1(32'hb689d4c4),
	.w2(32'hb932b37d),
	.w3(32'hb95624ec),
	.w4(32'hb8e241ab),
	.w5(32'hb9ae2fa8),
	.w6(32'h393de375),
	.w7(32'h3853ae94),
	.w8(32'hb950018c),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396ebc48),
	.w1(32'hb9a29db2),
	.w2(32'hb95b2c51),
	.w3(32'hba3918b8),
	.w4(32'hba96e8cc),
	.w5(32'hba9e6bb9),
	.w6(32'hba1d14c9),
	.w7(32'hba8510bf),
	.w8(32'hba847a60),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c2b233),
	.w1(32'hb9a1c637),
	.w2(32'hb950de16),
	.w3(32'h39155119),
	.w4(32'hba017fd0),
	.w5(32'hb8ffde24),
	.w6(32'h39aa8840),
	.w7(32'h386e67dd),
	.w8(32'h39b62ab9),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb983b2c5),
	.w1(32'hb917b111),
	.w2(32'hb7416dda),
	.w3(32'hb9991e81),
	.w4(32'h389c5ee3),
	.w5(32'h3910d5bf),
	.w6(32'hb9afc4fb),
	.w7(32'hb6ee3edc),
	.w8(32'h387f65d6),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a83eced),
	.w1(32'hb9a506f8),
	.w2(32'h3b029d81),
	.w3(32'hbac88c4f),
	.w4(32'hbad6085c),
	.w5(32'h3afa22fe),
	.w6(32'hbb1263e7),
	.w7(32'hbb29238e),
	.w8(32'h3a52309f),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a83ca31),
	.w1(32'h3ab1534c),
	.w2(32'h3a849436),
	.w3(32'hb9de6fa5),
	.w4(32'hba4be0d7),
	.w5(32'hbab63c8e),
	.w6(32'h3a1835e2),
	.w7(32'hb85f3b3d),
	.w8(32'hbad246e3),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388eabbc),
	.w1(32'hb6e305a8),
	.w2(32'h39a6348a),
	.w3(32'hb9adc920),
	.w4(32'hb9add935),
	.w5(32'h39416714),
	.w6(32'hb9107bda),
	.w7(32'h38dba3db),
	.w8(32'h38e31d3d),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h382ab386),
	.w1(32'h37b43fc8),
	.w2(32'h37b0dcd4),
	.w3(32'h37a9b4f0),
	.w4(32'h36ffe2d1),
	.w5(32'hb57a1d3d),
	.w6(32'hb78c8a62),
	.w7(32'h3719b6a3),
	.w8(32'hb8446176),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392cdab3),
	.w1(32'h3957c1a9),
	.w2(32'hb96a84f9),
	.w3(32'h380a12a2),
	.w4(32'hb8debb4f),
	.w5(32'hb9f27a5e),
	.w6(32'hb9a3e9f8),
	.w7(32'hba1a31bb),
	.w8(32'hba4dc422),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb829d236),
	.w1(32'hb80e2bd2),
	.w2(32'hb7f9f5ba),
	.w3(32'hb6fcbf8a),
	.w4(32'hb7bb3b8a),
	.w5(32'hb755a7d3),
	.w6(32'hb79fbbd6),
	.w7(32'hb7951538),
	.w8(32'h35ce26a1),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a53b273),
	.w1(32'h39ac4089),
	.w2(32'hb7a2e6cf),
	.w3(32'h39a22034),
	.w4(32'h3955fb5e),
	.w5(32'hb8fe4886),
	.w6(32'h38ac6fc2),
	.w7(32'hb997c7d0),
	.w8(32'hb9e79646),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94742cb),
	.w1(32'hb9b6e64e),
	.w2(32'hba08379f),
	.w3(32'hb8e298eb),
	.w4(32'hb9ce5933),
	.w5(32'hba51dc7e),
	.w6(32'h37f15e08),
	.w7(32'hb7afdfdd),
	.w8(32'hba596bd7),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d07b63),
	.w1(32'hb99e0839),
	.w2(32'hb9a612ca),
	.w3(32'hb9a78b93),
	.w4(32'hba54681b),
	.w5(32'hba6386e9),
	.w6(32'hba715d3a),
	.w7(32'hbaa663f7),
	.w8(32'hba9ae58e),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb81b1ff1),
	.w1(32'hb882de61),
	.w2(32'hb9d662d7),
	.w3(32'h391cae25),
	.w4(32'hb8bc25b6),
	.w5(32'hb9c7238f),
	.w6(32'hb9840061),
	.w7(32'hb9890d69),
	.w8(32'hb9a5e6de),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a219313),
	.w1(32'hba1bdfbf),
	.w2(32'h398bcf58),
	.w3(32'hba10a948),
	.w4(32'hbabeebbf),
	.w5(32'hb9a410c0),
	.w6(32'hba32828c),
	.w7(32'hbac8f17a),
	.w8(32'hba379038),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb921b2b6),
	.w1(32'h379731dd),
	.w2(32'h3976173f),
	.w3(32'hb9144189),
	.w4(32'hb915ab50),
	.w5(32'h39b779c1),
	.w6(32'hb7bd4113),
	.w7(32'h391b835d),
	.w8(32'h3a17bc7a),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h370de257),
	.w1(32'h3726753e),
	.w2(32'hb7653e44),
	.w3(32'h37c9dfc8),
	.w4(32'h37b67a02),
	.w5(32'hb6faf74b),
	.w6(32'h38090932),
	.w7(32'h373f5d3b),
	.w8(32'h36a0c00f),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a05a9c7),
	.w1(32'h39bda648),
	.w2(32'h3999fe6d),
	.w3(32'h39191d82),
	.w4(32'h382f552c),
	.w5(32'h39254a0a),
	.w6(32'h38cefd88),
	.w7(32'hb8da30f2),
	.w8(32'hb75eeb4f),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7f62ecb),
	.w1(32'h36aec92a),
	.w2(32'hb7dd9378),
	.w3(32'hb764dc6e),
	.w4(32'h37802175),
	.w5(32'hb6f69d5a),
	.w6(32'h3748b811),
	.w7(32'h3717f313),
	.w8(32'h37b83743),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a227542),
	.w1(32'h38d62635),
	.w2(32'h39843f03),
	.w3(32'hb90f96be),
	.w4(32'hba1e1847),
	.w5(32'hb97d4a8c),
	.w6(32'hb8fb65af),
	.w7(32'hba2b7c79),
	.w8(32'hb9d2a7b4),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3953f7fb),
	.w1(32'h3a56bbdd),
	.w2(32'h39118435),
	.w3(32'hba370206),
	.w4(32'h398888d4),
	.w5(32'hba6112b5),
	.w6(32'hb9c7016f),
	.w7(32'h3972c10b),
	.w8(32'hba1bff7c),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2278b3),
	.w1(32'h39008f45),
	.w2(32'h38f7556e),
	.w3(32'h3995aca0),
	.w4(32'hb9da5e82),
	.w5(32'hb974fc10),
	.w6(32'h38fc68ec),
	.w7(32'hba2a5c8e),
	.w8(32'hb9e5372d),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a11b49),
	.w1(32'hb933eba1),
	.w2(32'hb8dd890d),
	.w3(32'hb8d9cbeb),
	.w4(32'hb8929732),
	.w5(32'hb935561b),
	.w6(32'hb8c4914b),
	.w7(32'h388af909),
	.w8(32'hb94deb1f),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a74e8db),
	.w1(32'h37bb6d4b),
	.w2(32'hb977f62d),
	.w3(32'h39afae1f),
	.w4(32'hb9fc03f8),
	.w5(32'hb9f30fe0),
	.w6(32'hb8c4e3b6),
	.w7(32'hba6f2080),
	.w8(32'hba665639),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8f9596),
	.w1(32'hb93b2075),
	.w2(32'h39327dce),
	.w3(32'h3806dbff),
	.w4(32'hba901ecf),
	.w5(32'h3957c578),
	.w6(32'hba4b5520),
	.w7(32'hbade8a1c),
	.w8(32'hba1cf21b),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e4ba80),
	.w1(32'h3934f866),
	.w2(32'h394e3977),
	.w3(32'h39e37543),
	.w4(32'h3a1933b7),
	.w5(32'h39fb5f79),
	.w6(32'h39d3dc14),
	.w7(32'h3a18b6c3),
	.w8(32'h39d77fe3),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c4064e),
	.w1(32'hb7ddfa78),
	.w2(32'hb85f449b),
	.w3(32'hb8d66814),
	.w4(32'hb7cb3b54),
	.w5(32'hb836f335),
	.w6(32'hb87a4d2b),
	.w7(32'hb7e9aa95),
	.w8(32'hb844fa39),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb82514a1),
	.w1(32'h36206797),
	.w2(32'hb77c151a),
	.w3(32'hb7b6fb65),
	.w4(32'h36907bb1),
	.w5(32'hb6bae484),
	.w6(32'h361ee452),
	.w7(32'hb70cfa5c),
	.w8(32'hb31edcac),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0cc2dd),
	.w1(32'h3a1ec9b1),
	.w2(32'h3a142865),
	.w3(32'hba3ae84c),
	.w4(32'hb9d533fc),
	.w5(32'hba1f3ca1),
	.w6(32'hba5cae5a),
	.w7(32'hb9d2d0eb),
	.w8(32'hba2b43a8),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b110082),
	.w1(32'h3a564a4a),
	.w2(32'h39cf03f3),
	.w3(32'h3aa26778),
	.w4(32'hba7c0269),
	.w5(32'hb8c20a3c),
	.w6(32'h3a0b7531),
	.w7(32'hbadb8827),
	.w8(32'hb96d9a0c),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fa79e5),
	.w1(32'hb9bc3c42),
	.w2(32'hb92ae41b),
	.w3(32'hb8e4d97a),
	.w4(32'hba407d16),
	.w5(32'hb994628e),
	.w6(32'hb906084c),
	.w7(32'hba7c4de8),
	.w8(32'hba33a46a),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d5438c),
	.w1(32'h3a3763f9),
	.w2(32'h3a5bc76b),
	.w3(32'hba1525b0),
	.w4(32'hb9def195),
	.w5(32'h39e2e2d6),
	.w6(32'hba4318df),
	.w7(32'hb96094ed),
	.w8(32'hb95c54e2),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h380c8009),
	.w1(32'h37e916ca),
	.w2(32'h370889f3),
	.w3(32'hb76c7551),
	.w4(32'hb7d07b2d),
	.w5(32'hb8835194),
	.w6(32'h380ae268),
	.w7(32'hb886ee51),
	.w8(32'hb8615c4e),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0cc3a5),
	.w1(32'h39ef812a),
	.w2(32'h3934e6c8),
	.w3(32'h39cdcad9),
	.w4(32'h3981265b),
	.w5(32'h39508ed7),
	.w6(32'h395d10e1),
	.w7(32'h3921b164),
	.w8(32'h3997bc26),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7e79dc8),
	.w1(32'hb9a8d031),
	.w2(32'h389ad97c),
	.w3(32'h381d550c),
	.w4(32'h389c27a3),
	.w5(32'h38a28868),
	.w6(32'h3a4bba03),
	.w7(32'h38b299a5),
	.w8(32'hb72c6344),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8dd9b1),
	.w1(32'h3a798306),
	.w2(32'h3abc82ad),
	.w3(32'hb814f3ff),
	.w4(32'h39995e95),
	.w5(32'h39f2138e),
	.w6(32'hb84ca58e),
	.w7(32'h3958b68e),
	.w8(32'h3a28e4e1),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1e6987),
	.w1(32'h38defc90),
	.w2(32'h39ccadb0),
	.w3(32'hb94a9a61),
	.w4(32'hba20c730),
	.w5(32'hb90da8fd),
	.w6(32'h38b62304),
	.w7(32'hb9d2797a),
	.w8(32'hb7526f3c),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397d4eb0),
	.w1(32'h39e70f98),
	.w2(32'hb9936f14),
	.w3(32'hb917188d),
	.w4(32'h38f0201f),
	.w5(32'hba79e90b),
	.w6(32'h391b7020),
	.w7(32'h39d46159),
	.w8(32'hba520fd8),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a896e09),
	.w1(32'h3a0a96c9),
	.w2(32'hb9abaeeb),
	.w3(32'h39ad2156),
	.w4(32'hb982848e),
	.w5(32'hba8cb8ff),
	.w6(32'hb8964b6b),
	.w7(32'hba4b510c),
	.w8(32'hbaa23ea5),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7d87256),
	.w1(32'hb734a307),
	.w2(32'hb74a03a3),
	.w3(32'hb7b5fd02),
	.w4(32'hb4ff5262),
	.w5(32'hb7025e6f),
	.w6(32'hb58e7a1a),
	.w7(32'h36f0b9f7),
	.w8(32'hb728ae28),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb73c3884),
	.w1(32'hb5ef111f),
	.w2(32'hb76c5336),
	.w3(32'hb6c2ff68),
	.w4(32'hb6a7801c),
	.w5(32'hb7a9d201),
	.w6(32'hb704fadf),
	.w7(32'hb6c3741d),
	.w8(32'h3631014a),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37e84812),
	.w1(32'h38a48cae),
	.w2(32'h389b3cf8),
	.w3(32'hb9d523ba),
	.w4(32'h38051bfe),
	.w5(32'hb751dfb1),
	.w6(32'hb92b1eb0),
	.w7(32'hb88043ad),
	.w8(32'h383d594f),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb60f081f),
	.w1(32'h36b0e741),
	.w2(32'hb65fd4f3),
	.w3(32'h374c2d46),
	.w4(32'h3802f305),
	.w5(32'h35901312),
	.w6(32'h37ecfa49),
	.w7(32'h379274cd),
	.w8(32'hb783a935),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8938b4b),
	.w1(32'h393d97ff),
	.w2(32'h396f5c52),
	.w3(32'hb8e27bab),
	.w4(32'h39c64899),
	.w5(32'h39babe58),
	.w6(32'hb8d4efd1),
	.w7(32'h39afe7eb),
	.w8(32'h393433b3),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aca72cf),
	.w1(32'hb886bd56),
	.w2(32'hb8639f97),
	.w3(32'h3a47fd83),
	.w4(32'hba415c0c),
	.w5(32'hb9b25060),
	.w6(32'h3996ebaa),
	.w7(32'hbaa3bef3),
	.w8(32'hba92defd),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399c1ea0),
	.w1(32'hb9c49048),
	.w2(32'hb907177b),
	.w3(32'h39c0ff07),
	.w4(32'hb9ab0c0e),
	.w5(32'h35acf360),
	.w6(32'h3868c9ed),
	.w7(32'hba667c45),
	.w8(32'hba003255),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37be02b4),
	.w1(32'h374b20e7),
	.w2(32'hb786b412),
	.w3(32'h37b7d02c),
	.w4(32'hb6dddf17),
	.w5(32'hb7ec292d),
	.w6(32'h34bc5a0d),
	.w7(32'h37541905),
	.w8(32'h371449bf),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac9e352),
	.w1(32'h39956b49),
	.w2(32'h3a3cd9fd),
	.w3(32'hb970755b),
	.w4(32'hba7d33db),
	.w5(32'hb9112798),
	.w6(32'hb992bfc6),
	.w7(32'hba683aeb),
	.w8(32'hb879f9d2),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a510f9c),
	.w1(32'h3946f27b),
	.w2(32'h39eecfc5),
	.w3(32'hb94b9fcb),
	.w4(32'hb9d46ecb),
	.w5(32'h37cbe4c0),
	.w6(32'hb9c90168),
	.w7(32'hb9da0e19),
	.w8(32'h3926272c),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38418aab),
	.w1(32'hb9b0b0d5),
	.w2(32'hb91cf3e4),
	.w3(32'hb917ab1f),
	.w4(32'hba04c406),
	.w5(32'hb9daaa1a),
	.w6(32'hb973e362),
	.w7(32'hb9fc90ea),
	.w8(32'hb99eed35),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39caf813),
	.w1(32'h397f6f53),
	.w2(32'h3a246dbc),
	.w3(32'hb97eb184),
	.w4(32'hb9479f19),
	.w5(32'h39bfbccb),
	.w6(32'hb95a5d5e),
	.w7(32'hb98b213c),
	.w8(32'h38888a67),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7b4448a),
	.w1(32'hb9279eda),
	.w2(32'hb963debc),
	.w3(32'hb8e7bf42),
	.w4(32'hb93ccd77),
	.w5(32'hb92a9d42),
	.w6(32'hb932344b),
	.w7(32'hb97e1946),
	.w8(32'hb9282084),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3762eec1),
	.w1(32'h3869323d),
	.w2(32'h3893a740),
	.w3(32'h3887e645),
	.w4(32'h39102bd7),
	.w5(32'h38c50a95),
	.w6(32'h37b02a5d),
	.w7(32'h36ec400b),
	.w8(32'h3706c4ce),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h362853c4),
	.w1(32'h37f2adab),
	.w2(32'h37a58c6c),
	.w3(32'hb7f5c99c),
	.w4(32'hb7330615),
	.w5(32'hb766bb3e),
	.w6(32'hb7a3401d),
	.w7(32'hb7ffc17c),
	.w8(32'h372fa2ae),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88e845e),
	.w1(32'hb806b5d1),
	.w2(32'hb786b7a7),
	.w3(32'hb83d57a9),
	.w4(32'hb72f66b0),
	.w5(32'h367c51eb),
	.w6(32'hb8434029),
	.w7(32'h371821bf),
	.w8(32'hb79e1663),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d5806a),
	.w1(32'h38a71e41),
	.w2(32'hba373d07),
	.w3(32'hb9670ac2),
	.w4(32'hb942aa08),
	.w5(32'hba8856af),
	.w6(32'h391e920a),
	.w7(32'h38ef8e17),
	.w8(32'hba96fec5),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a537e14),
	.w1(32'hb9832dd0),
	.w2(32'h3a563b70),
	.w3(32'hb817a14e),
	.w4(32'hba93fb1a),
	.w5(32'h3a3683f9),
	.w6(32'hba4a2f13),
	.w7(32'hbae7d439),
	.w8(32'hb9c2377a),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af2efda),
	.w1(32'h3a403e50),
	.w2(32'h3a850a31),
	.w3(32'h39f28514),
	.w4(32'hba5afd18),
	.w5(32'h38718855),
	.w6(32'hba361548),
	.w7(32'hbadcd745),
	.w8(32'hba280393),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a17f4d6),
	.w1(32'hb805b045),
	.w2(32'h3a381153),
	.w3(32'hb93f4a94),
	.w4(32'hba32a453),
	.w5(32'h3a39e2ab),
	.w6(32'h3947fe63),
	.w7(32'hba0d548f),
	.w8(32'h396c3b51),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a3e4cc),
	.w1(32'hb904d1e4),
	.w2(32'hb948d099),
	.w3(32'hb8e454d5),
	.w4(32'hb918efdd),
	.w5(32'hb947c6ae),
	.w6(32'hb849d001),
	.w7(32'hb8b15815),
	.w8(32'hb934b07a),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e036c9),
	.w1(32'h3797ca2b),
	.w2(32'h371348f9),
	.w3(32'hb7bd9e59),
	.w4(32'h3811fccb),
	.w5(32'h379d9017),
	.w6(32'hb8784ab6),
	.w7(32'hb89f2c4b),
	.w8(32'h36c8f6ce),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38bd9327),
	.w1(32'h39121d83),
	.w2(32'h36755741),
	.w3(32'h383ac979),
	.w4(32'h388e741e),
	.w5(32'h38467a94),
	.w6(32'h38567f29),
	.w7(32'h3873336f),
	.w8(32'h38672059),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5350276),
	.w1(32'h37614855),
	.w2(32'h37955da6),
	.w3(32'hb8348245),
	.w4(32'hb7c7f9b6),
	.w5(32'hb7e9754b),
	.w6(32'hb8137c22),
	.w7(32'hb8790658),
	.w8(32'hb84402dd),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4a83d5),
	.w1(32'h39a06501),
	.w2(32'h3a0e0fe7),
	.w3(32'h39e87de7),
	.w4(32'hb88880a8),
	.w5(32'hb8c89a57),
	.w6(32'hb8b591e2),
	.w7(32'hb9483f94),
	.w8(32'h37a0ce80),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a181fe),
	.w1(32'h38442e1a),
	.w2(32'hb912c972),
	.w3(32'h39836095),
	.w4(32'hb7a28e93),
	.w5(32'hb96715fb),
	.w6(32'hb64c3369),
	.w7(32'hb9957b96),
	.w8(32'hb9a0c018),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2cf62b),
	.w1(32'hb915912c),
	.w2(32'hb990e334),
	.w3(32'hba281a40),
	.w4(32'hb907d8be),
	.w5(32'hb9a5a5df),
	.w6(32'hba0645da),
	.w7(32'hb854c31b),
	.w8(32'hb9c51a50),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92785fd),
	.w1(32'hb84bc232),
	.w2(32'hb854e227),
	.w3(32'hb8d99fd6),
	.w4(32'hb8a999ef),
	.w5(32'hb899f017),
	.w6(32'hb7dccec0),
	.w7(32'h367a2e9d),
	.w8(32'h3838c90f),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38df2995),
	.w1(32'h380d6e2c),
	.w2(32'hb8cca961),
	.w3(32'h37af47e4),
	.w4(32'hb8cea05c),
	.w5(32'hb8e7fdfb),
	.w6(32'h3866a2f1),
	.w7(32'hb971cc70),
	.w8(32'hb90d5ef5),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393eecda),
	.w1(32'h393c14c6),
	.w2(32'h39569a71),
	.w3(32'hb8475093),
	.w4(32'h3793c51b),
	.w5(32'h37e4796b),
	.w6(32'h368590dd),
	.w7(32'hb7d528fe),
	.w8(32'h38687ae8),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37154a5b),
	.w1(32'h38046e56),
	.w2(32'hb83c78eb),
	.w3(32'hb867e073),
	.w4(32'h37842e6a),
	.w5(32'hb83c07e3),
	.w6(32'hb8db8a1d),
	.w7(32'hb85bea39),
	.w8(32'hb83809cc),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb841e0c6),
	.w1(32'h3945ce36),
	.w2(32'h3a8c1429),
	.w3(32'hb9936d93),
	.w4(32'hb9fe7395),
	.w5(32'hb8de7586),
	.w6(32'hbade9c94),
	.w7(32'hbabbd74d),
	.w8(32'hba4480f6),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6e41aae),
	.w1(32'hbb838585),
	.w2(32'hb9e4b600),
	.w3(32'hb7b81cbf),
	.w4(32'h39ce8b21),
	.w5(32'h3ba3d1b3),
	.w6(32'hbb709b78),
	.w7(32'hbb5c91a6),
	.w8(32'h3ab0a5e3),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5be39d),
	.w1(32'h3b44d24f),
	.w2(32'h3bceded8),
	.w3(32'h3a0ec9c5),
	.w4(32'hbaaa4928),
	.w5(32'h3a69af5c),
	.w6(32'hbb5c175f),
	.w7(32'hba669e2b),
	.w8(32'h3adeb5f4),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule