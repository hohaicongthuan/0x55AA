module layer_6_featuremap_90(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 2048;
	parameter IMG_SIZE = 52;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbcd902),
	.w1(32'hbb3595a6),
	.w2(32'h3b0697a7),
	.w3(32'h3b8f5155),
	.w4(32'hbb6c107b),
	.w5(32'hbaf1be93),
	.w6(32'h3af79531),
	.w7(32'hbaa7978c),
	.w8(32'h3a532591),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3c9db2),
	.w1(32'h3b17b0ed),
	.w2(32'h3c0529fb),
	.w3(32'hb905f3de),
	.w4(32'h3afc2ab3),
	.w5(32'h3ab70e9b),
	.w6(32'h3b21ecec),
	.w7(32'hb9decf4e),
	.w8(32'h3a12bc0c),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba83607),
	.w1(32'h3cd07be0),
	.w2(32'h3a2aaf0f),
	.w3(32'hbd15efe8),
	.w4(32'h3ce66d65),
	.w5(32'hbb3211dd),
	.w6(32'h3b9a63c5),
	.w7(32'h3ca4cadb),
	.w8(32'hbc816e7a),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc69f101),
	.w1(32'h3b2da889),
	.w2(32'h3ab4df45),
	.w3(32'hba242438),
	.w4(32'h3b476076),
	.w5(32'h3b0df548),
	.w6(32'h396db9d9),
	.w7(32'h3b90cf3c),
	.w8(32'hbab08b49),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6a6666),
	.w1(32'hbcf45473),
	.w2(32'h3cd2e17e),
	.w3(32'h3c13230a),
	.w4(32'hbd036f73),
	.w5(32'h3be2900b),
	.w6(32'hbbf16b00),
	.w7(32'hbd2e4307),
	.w8(32'h3cc38796),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaf7a49),
	.w1(32'hbb701f6f),
	.w2(32'hbb04045d),
	.w3(32'h3bb0d5a0),
	.w4(32'hba9c0a6d),
	.w5(32'hbb50d16d),
	.w6(32'h3a0218b0),
	.w7(32'hbb21f4f0),
	.w8(32'hbb81e4ef),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb92c8ad),
	.w1(32'hbb4084c5),
	.w2(32'hbbcd5cb1),
	.w3(32'hbb84e0ed),
	.w4(32'h3b39e003),
	.w5(32'hbb29fba3),
	.w6(32'hbb1c3d14),
	.w7(32'hbac0bd78),
	.w8(32'h3b885e93),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b444084),
	.w1(32'hbb947525),
	.w2(32'hbd2c1764),
	.w3(32'hbb97b283),
	.w4(32'h3ca06315),
	.w5(32'hbc7e2d69),
	.w6(32'h3c5ad04b),
	.w7(32'hbcab30d6),
	.w8(32'hbcca8066),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c86eab4),
	.w1(32'h3ca785e8),
	.w2(32'h3c591e6b),
	.w3(32'hbc908c59),
	.w4(32'h3b1382db),
	.w5(32'h3c83127b),
	.w6(32'hbcac984a),
	.w7(32'h3d4b4519),
	.w8(32'hbcec9b85),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbaa139),
	.w1(32'h3a9fe006),
	.w2(32'h3bc3a089),
	.w3(32'h3b897875),
	.w4(32'hba9136c0),
	.w5(32'h3b53c877),
	.w6(32'h39e25d37),
	.w7(32'h3bb20a0a),
	.w8(32'hb933fb2d),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab70428),
	.w1(32'h3c1435b3),
	.w2(32'h3d4fb3e7),
	.w3(32'h3c977adc),
	.w4(32'h3bf7e5b2),
	.w5(32'h3cfd653f),
	.w6(32'h3cf6ccdd),
	.w7(32'h3d43eb12),
	.w8(32'h3d3ce729),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba48a318),
	.w1(32'h3a3a6f83),
	.w2(32'h3c2bcc3d),
	.w3(32'h3c38cac8),
	.w4(32'hbbad33fe),
	.w5(32'h3a953636),
	.w6(32'hbb42da15),
	.w7(32'hbb0b0dea),
	.w8(32'hbb0fc5f5),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc08e7dc),
	.w1(32'hbb752b68),
	.w2(32'h3c71335e),
	.w3(32'h3abdcf58),
	.w4(32'h3c58f149),
	.w5(32'hbb767602),
	.w6(32'hba3f3bbe),
	.w7(32'h3c9c5be0),
	.w8(32'hbb81c0d4),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7cfad8),
	.w1(32'h3b91544f),
	.w2(32'h3b867d4f),
	.w3(32'hbbb43ddd),
	.w4(32'hbc1aedfe),
	.w5(32'hbb021d56),
	.w6(32'hbbaa912f),
	.w7(32'hbb82f96c),
	.w8(32'h3b80fc69),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b770595),
	.w1(32'h3b0b3a26),
	.w2(32'h3bf35d53),
	.w3(32'hb8bf708a),
	.w4(32'hba14318f),
	.w5(32'hbb8232da),
	.w6(32'hbaadf6e5),
	.w7(32'h3b508445),
	.w8(32'h3ad1a5f8),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2990d5),
	.w1(32'h3b2d6de7),
	.w2(32'hba1a0eaf),
	.w3(32'hbb00be94),
	.w4(32'h3a7f77eb),
	.w5(32'hbbad89b8),
	.w6(32'h398aeed0),
	.w7(32'h393fe542),
	.w8(32'hbb8febc2),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c01a802),
	.w1(32'h3cb4f3dd),
	.w2(32'h3c033dcf),
	.w3(32'h3bf2bd65),
	.w4(32'h3cb6d8d5),
	.w5(32'h3b03d235),
	.w6(32'h3c0e4614),
	.w7(32'h3ca7082a),
	.w8(32'hbc37cafb),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6925e5),
	.w1(32'hbb5f256c),
	.w2(32'hbbc7c3ce),
	.w3(32'h3b9ab6fa),
	.w4(32'hba1824ea),
	.w5(32'h3a430024),
	.w6(32'hba43364d),
	.w7(32'hba18567e),
	.w8(32'hbb49e674),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1f8ea9),
	.w1(32'h3a80580f),
	.w2(32'hb8b71cb1),
	.w3(32'h399f8f19),
	.w4(32'h38c0c856),
	.w5(32'h39293368),
	.w6(32'h3b03c8d4),
	.w7(32'hba0b93be),
	.w8(32'h3a0cbd67),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab062b9),
	.w1(32'hbbcbdc33),
	.w2(32'h3b75b0d7),
	.w3(32'h3b328734),
	.w4(32'hbc7a0c19),
	.w5(32'hbcf73989),
	.w6(32'h3c0b98fc),
	.w7(32'hbcc2fb86),
	.w8(32'hbc20c1c4),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc57e1fb),
	.w1(32'hba3ebc66),
	.w2(32'hbaaaf365),
	.w3(32'hbb2574d3),
	.w4(32'h3ac90d89),
	.w5(32'hba1a953a),
	.w6(32'hbb3909f3),
	.w7(32'hb7fc956e),
	.w8(32'h3a30d6a7),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1ccd8f),
	.w1(32'h3be33ea2),
	.w2(32'h3c760004),
	.w3(32'hbb0ab8ef),
	.w4(32'h3b232d89),
	.w5(32'h3b261a30),
	.w6(32'h3b35177f),
	.w7(32'h3c44be5e),
	.w8(32'h3b69fc67),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7c520b),
	.w1(32'h3b1f0e94),
	.w2(32'h3be52a5b),
	.w3(32'hbbcf180a),
	.w4(32'hbb314800),
	.w5(32'h3c6db797),
	.w6(32'hbce77b9e),
	.w7(32'h3cc86d77),
	.w8(32'hbc9847f4),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb203e2),
	.w1(32'h3c853645),
	.w2(32'hbaf85f30),
	.w3(32'hba0820e1),
	.w4(32'h3d07133a),
	.w5(32'hbc90b82c),
	.w6(32'h3c0796e3),
	.w7(32'h3bbcf5b1),
	.w8(32'hbc85cabe),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba5fbeb),
	.w1(32'h3c7e44e1),
	.w2(32'h398a41b6),
	.w3(32'hbc88de37),
	.w4(32'h3bdbb069),
	.w5(32'hbc3d756d),
	.w6(32'h3bc482bf),
	.w7(32'h3c19fcc2),
	.w8(32'hbc221a4f),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b99cd44),
	.w1(32'h3b9671c6),
	.w2(32'hbb03ba10),
	.w3(32'hb9fc0991),
	.w4(32'h3c094a19),
	.w5(32'h3b28916e),
	.w6(32'h3bd80578),
	.w7(32'hba3fdbb0),
	.w8(32'hba815164),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3ea1ec),
	.w1(32'h3b8d5538),
	.w2(32'h3c4a4c81),
	.w3(32'h38f2f705),
	.w4(32'h3b973533),
	.w5(32'h3b6f361e),
	.w6(32'h3b386222),
	.w7(32'h3c77479c),
	.w8(32'h3b6ef55e),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7c79b9),
	.w1(32'h3b0ac54d),
	.w2(32'hbb2cdf84),
	.w3(32'hbbf5927a),
	.w4(32'h3b5bd9e5),
	.w5(32'hbac647df),
	.w6(32'h39ef7443),
	.w7(32'hbb864ac5),
	.w8(32'h3b415e6b),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb167c6),
	.w1(32'h3b2669a7),
	.w2(32'h3b27d1e4),
	.w3(32'hbba5cd5a),
	.w4(32'hb9d4c627),
	.w5(32'hbaa091bf),
	.w6(32'h3ad76fe4),
	.w7(32'h3ac6b8d4),
	.w8(32'h3b1afb16),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbeb993),
	.w1(32'hbd02c8c6),
	.w2(32'h3c440f73),
	.w3(32'h3c29ae3c),
	.w4(32'h3c86ae8b),
	.w5(32'h3bbf9441),
	.w6(32'hbccca9f6),
	.w7(32'h3c350775),
	.w8(32'h3cd62b42),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc26f0ba),
	.w1(32'h3ca90046),
	.w2(32'hbd10f000),
	.w3(32'h3a856983),
	.w4(32'h3cb7a73f),
	.w5(32'hbd329307),
	.w6(32'h3ca0f028),
	.w7(32'hbcbe3fe7),
	.w8(32'h3ae5257c),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cf8d2c4),
	.w1(32'hbc1f8058),
	.w2(32'h3bc3c20c),
	.w3(32'h3ca5578c),
	.w4(32'hbbe585f6),
	.w5(32'h3ae01187),
	.w6(32'h3c0224ed),
	.w7(32'hbc13bf48),
	.w8(32'h3b125ef4),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba34e99f),
	.w1(32'h3c76ed77),
	.w2(32'hbca6918e),
	.w3(32'h3a78a637),
	.w4(32'h3ca47e46),
	.w5(32'hbc98000b),
	.w6(32'hbb5023a2),
	.w7(32'h3c8aafc0),
	.w8(32'hbd03ac19),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a434da3),
	.w1(32'h3aef374b),
	.w2(32'h38406e6d),
	.w3(32'hbbd9b4b6),
	.w4(32'h3c18fa4f),
	.w5(32'hbbb81e74),
	.w6(32'hbc10ce5b),
	.w7(32'hbafae75a),
	.w8(32'hbbc86148),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b93d968),
	.w1(32'hbb66e769),
	.w2(32'h3b8013da),
	.w3(32'h3af1e747),
	.w4(32'hbabb74e7),
	.w5(32'hba827be5),
	.w6(32'hba914fdf),
	.w7(32'h3b22ef2c),
	.w8(32'hbb60b9a7),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc1306c),
	.w1(32'hbb5bca3d),
	.w2(32'h3c648914),
	.w3(32'h3bf8ccfc),
	.w4(32'h3c030e1c),
	.w5(32'h3c4af010),
	.w6(32'hbbd7def5),
	.w7(32'h3b9c5a5b),
	.w8(32'h3bbae9fb),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4cd15b),
	.w1(32'hb95af30e),
	.w2(32'h3b4b4133),
	.w3(32'h3b6c5b17),
	.w4(32'hb9a18136),
	.w5(32'h3a6af05c),
	.w6(32'h3b7f4971),
	.w7(32'hbbe6c151),
	.w8(32'hba3042fc),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc34f6c3),
	.w1(32'h39050939),
	.w2(32'hba3236ff),
	.w3(32'hbb63b0dc),
	.w4(32'h3abbee63),
	.w5(32'hbb2c9b0f),
	.w6(32'hb9c8fcfd),
	.w7(32'hbb842d9c),
	.w8(32'hb8b28317),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b299bac),
	.w1(32'hbc51d17f),
	.w2(32'hbc268f12),
	.w3(32'hbcb0d767),
	.w4(32'hbc65d755),
	.w5(32'hbc47155d),
	.w6(32'hbbfa93af),
	.w7(32'hbc9ddd8c),
	.w8(32'hbc87b3b5),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba03610),
	.w1(32'hbcdfec08),
	.w2(32'hbcd96087),
	.w3(32'h3cb80fa7),
	.w4(32'h3c30f589),
	.w5(32'hbd5f4d81),
	.w6(32'h3cfa85a2),
	.w7(32'hbda85d4e),
	.w8(32'h3d166ed9),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cccfa21),
	.w1(32'h3ccc1252),
	.w2(32'hbc5a6efe),
	.w3(32'h3c962264),
	.w4(32'h3c7cfa8e),
	.w5(32'hbd4148e3),
	.w6(32'h3d227657),
	.w7(32'hbcd0edae),
	.w8(32'h3bea421d),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb1b6c2),
	.w1(32'h3b68c500),
	.w2(32'h3ba9c82a),
	.w3(32'hba8d62a2),
	.w4(32'h3bab0f94),
	.w5(32'h3b1c5b32),
	.w6(32'hb7bb2340),
	.w7(32'h3ba6407e),
	.w8(32'h3b3a0e20),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8ef29b),
	.w1(32'h3c13172f),
	.w2(32'h3b6e60fb),
	.w3(32'h3c068e1f),
	.w4(32'h3b419033),
	.w5(32'h3b84efad),
	.w6(32'h3c0a54d4),
	.w7(32'h3be4e688),
	.w8(32'hb8efa388),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce41b20),
	.w1(32'hbcb5b04f),
	.w2(32'hbb6ce56c),
	.w3(32'h3bf16e05),
	.w4(32'h3cce8dbf),
	.w5(32'h3c3b9d9c),
	.w6(32'hbc1bc2bc),
	.w7(32'h3be9dd7d),
	.w8(32'h3bc5c5f5),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2be61b),
	.w1(32'h3c06ec8e),
	.w2(32'h3bbf8548),
	.w3(32'hbaacea2a),
	.w4(32'hba82d4f5),
	.w5(32'hbb9442ee),
	.w6(32'h3b762e62),
	.w7(32'h3ba1a9ba),
	.w8(32'h38cff862),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b46126),
	.w1(32'hbc1d8de5),
	.w2(32'h3cd6f455),
	.w3(32'h3c50562e),
	.w4(32'h3bb18ee1),
	.w5(32'h3bcf5b23),
	.w6(32'h3b745dd3),
	.w7(32'h3c7686ad),
	.w8(32'h3c987d69),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcdf9b93),
	.w1(32'h3af0bfdc),
	.w2(32'h3b29e1db),
	.w3(32'hbb20fc1f),
	.w4(32'h3c0ead9f),
	.w5(32'hbc4923c7),
	.w6(32'hba80f74b),
	.w7(32'h3ad67e44),
	.w8(32'hbc3d8937),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c17ce98),
	.w1(32'hbc53aa31),
	.w2(32'hbce4c9c6),
	.w3(32'hbbb5218a),
	.w4(32'hbcc8a12c),
	.w5(32'hbcf92a39),
	.w6(32'hbc7cee28),
	.w7(32'hbd1642f0),
	.w8(32'hbd28d9a1),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbccdae06),
	.w1(32'hba6893ef),
	.w2(32'h39ab6e1c),
	.w3(32'h3bd31513),
	.w4(32'h38b7b4e0),
	.w5(32'hbb7c631f),
	.w6(32'h3ac1285d),
	.w7(32'hbada102a),
	.w8(32'hbad09d6b),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb367fea),
	.w1(32'hbd0e3a33),
	.w2(32'hbc56a31f),
	.w3(32'h3ca63dae),
	.w4(32'hbc8e18ba),
	.w5(32'hbcbdaf08),
	.w6(32'h3c98d4dc),
	.w7(32'hbd6f6bb0),
	.w8(32'h3ce8a8ca),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d1375a3),
	.w1(32'h3b430aa1),
	.w2(32'h3bcc59b3),
	.w3(32'hb9f48634),
	.w4(32'h3c0e223d),
	.w5(32'h3acd0f40),
	.w6(32'hb8afdd7d),
	.w7(32'h3c336112),
	.w8(32'h3ab33d93),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6204c2),
	.w1(32'h3b9c37ec),
	.w2(32'h3b7ce6df),
	.w3(32'hb75d517a),
	.w4(32'h3be635bb),
	.w5(32'h3bc9aae9),
	.w6(32'h3b4c2f3c),
	.w7(32'h3af0f679),
	.w8(32'h3bd49178),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c543964),
	.w1(32'h3cbd717a),
	.w2(32'h3c091e7d),
	.w3(32'h3ba298bf),
	.w4(32'h3c1f0599),
	.w5(32'h38e5c8e3),
	.w6(32'h3ca02c52),
	.w7(32'h3c1714d4),
	.w8(32'hba174ccd),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2eede9),
	.w1(32'hbb3fb124),
	.w2(32'hbbf68153),
	.w3(32'hbb2047dc),
	.w4(32'hbb932da9),
	.w5(32'hbc5561e4),
	.w6(32'hbafd0aca),
	.w7(32'hbb98040a),
	.w8(32'hbc0e495b),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba25725),
	.w1(32'hbaaa7369),
	.w2(32'h3a9427bb),
	.w3(32'h3ab51d03),
	.w4(32'h3b7e66d7),
	.w5(32'h3a996891),
	.w6(32'h3ab5a53e),
	.w7(32'h3bc2438d),
	.w8(32'hba0d80fa),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f8ced3),
	.w1(32'hbb8b0805),
	.w2(32'hbb02e1fc),
	.w3(32'h3c48a765),
	.w4(32'h3ad185a6),
	.w5(32'hbb706e0e),
	.w6(32'hbcc855a8),
	.w7(32'hbd26934b),
	.w8(32'hbd059f3e),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c954aab),
	.w1(32'hbc1fa763),
	.w2(32'hbc3270e8),
	.w3(32'h3c4517bb),
	.w4(32'h3cb92856),
	.w5(32'h3c6b47a1),
	.w6(32'h3bc76553),
	.w7(32'h3c26ac7f),
	.w8(32'h3bfe3007),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc07f696),
	.w1(32'hbbabde24),
	.w2(32'h3b09c92a),
	.w3(32'hbbcd74e4),
	.w4(32'hbc8908ff),
	.w5(32'hbb2ae8b2),
	.w6(32'hbc175936),
	.w7(32'hbccad6db),
	.w8(32'hbbbfd3ca),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad7d3fe),
	.w1(32'h3b88c9fe),
	.w2(32'h3c092d93),
	.w3(32'hbc22f2a1),
	.w4(32'hbc406901),
	.w5(32'hbbd08637),
	.w6(32'hbb8c23fa),
	.w7(32'hbae858ee),
	.w8(32'h3b18cffb),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2fc371),
	.w1(32'h3c9d2e28),
	.w2(32'h3cc90949),
	.w3(32'hbba1e83d),
	.w4(32'hbcd12cda),
	.w5(32'hbcfff7b6),
	.w6(32'hbc1130e6),
	.w7(32'hbc20b70e),
	.w8(32'hba1c905c),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c720acd),
	.w1(32'h3c153118),
	.w2(32'h3c8aa735),
	.w3(32'hba280889),
	.w4(32'hbc24f8b1),
	.w5(32'hbc125c2d),
	.w6(32'h3b9d9bed),
	.w7(32'h3b88ab6d),
	.w8(32'h3b48f2ca),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca32f74),
	.w1(32'h3cbe41bf),
	.w2(32'h3ccf515b),
	.w3(32'h3c913c6e),
	.w4(32'h3ccdd06f),
	.w5(32'h3c33ff55),
	.w6(32'h3c9b7fce),
	.w7(32'h3caaa7e1),
	.w8(32'h3c9df2ef),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c698491),
	.w1(32'hbd276f3e),
	.w2(32'hbd378636),
	.w3(32'h3ceb54c2),
	.w4(32'h3d32a14c),
	.w5(32'h3c7b97c2),
	.w6(32'hbce75298),
	.w7(32'hbbef01f0),
	.w8(32'h3bdcfe0b),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1b4d89),
	.w1(32'h3c9f5ac2),
	.w2(32'h3d2b910e),
	.w3(32'hbd037d0b),
	.w4(32'hbd26322c),
	.w5(32'hbcfedf00),
	.w6(32'hbb98b637),
	.w7(32'h3b1b25e5),
	.w8(32'h3b6a7eab),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

endmodule