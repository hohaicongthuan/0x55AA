module layer_10_featuremap_95(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba221cda),
	.w1(32'h3b8d8f59),
	.w2(32'hb9facc1c),
	.w3(32'hb9c43075),
	.w4(32'h3b9ee64c),
	.w5(32'hba20f0b1),
	.w6(32'h3b6def38),
	.w7(32'hba58a3e1),
	.w8(32'h3a534a79),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2a029f),
	.w1(32'hbab3fb57),
	.w2(32'h3aa2d377),
	.w3(32'h3a887dcc),
	.w4(32'hba99fbd4),
	.w5(32'h3a85c28b),
	.w6(32'hb93da64e),
	.w7(32'h3a92f432),
	.w8(32'h39735be1),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1ad54b),
	.w1(32'hbaa21c90),
	.w2(32'hbaa59917),
	.w3(32'hb90227ba),
	.w4(32'hbae0bb9b),
	.w5(32'hbadebaac),
	.w6(32'hbab09d60),
	.w7(32'hbaceeb1e),
	.w8(32'hbb015af2),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeec301),
	.w1(32'hbb27ce59),
	.w2(32'hbb52a003),
	.w3(32'hbb113095),
	.w4(32'hba31a06a),
	.w5(32'hb99b8cd2),
	.w6(32'hbac7e0e4),
	.w7(32'hbb63dc31),
	.w8(32'hbb0bcd36),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1c386a),
	.w1(32'h3af97280),
	.w2(32'h3a1a8470),
	.w3(32'hba593215),
	.w4(32'h3ade1434),
	.w5(32'h3a26368b),
	.w6(32'h3b043009),
	.w7(32'h396f92d1),
	.w8(32'hbaddf059),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2cc74b),
	.w1(32'hbaa09e5c),
	.w2(32'hbaceae32),
	.w3(32'hba21dc52),
	.w4(32'hbad1eb15),
	.w5(32'hbb091bc1),
	.w6(32'hba2c3f98),
	.w7(32'hbabdd857),
	.w8(32'h39e17176),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a15eeef),
	.w1(32'hbaa4292f),
	.w2(32'h3a097f81),
	.w3(32'hb9f75309),
	.w4(32'hbaa3d0bb),
	.w5(32'h39cba43d),
	.w6(32'hba8f57fa),
	.w7(32'h3a4b8c19),
	.w8(32'hba388fc2),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa71fad),
	.w1(32'h39694395),
	.w2(32'hba96a248),
	.w3(32'hba8332c9),
	.w4(32'h3abe1f16),
	.w5(32'h38fdf72d),
	.w6(32'h3a4c33ec),
	.w7(32'hba8c0f30),
	.w8(32'h3918d84a),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb984dc55),
	.w1(32'h3b3d21cf),
	.w2(32'h39811181),
	.w3(32'h3a0378b6),
	.w4(32'h3b2f52c8),
	.w5(32'hb9a9257f),
	.w6(32'h3b300394),
	.w7(32'hb93995a4),
	.w8(32'hb89e886f),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba58fc87),
	.w1(32'hb9dd9922),
	.w2(32'h3a12c7f9),
	.w3(32'hb9a8ca18),
	.w4(32'h3a3634c1),
	.w5(32'h3aedb58f),
	.w6(32'h3a454a41),
	.w7(32'h3b080607),
	.w8(32'h3b469f4c),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acdc953),
	.w1(32'hbb1a6038),
	.w2(32'hba4bee81),
	.w3(32'h3afc0658),
	.w4(32'hbb8e0c1f),
	.w5(32'hbac70c11),
	.w6(32'hbb38b61a),
	.w7(32'hbb18d58e),
	.w8(32'hba30f090),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9467fbc),
	.w1(32'hb9f2e385),
	.w2(32'h3ab22c45),
	.w3(32'hb9fa8f40),
	.w4(32'hbac10b0c),
	.w5(32'hb6809f23),
	.w6(32'hba65405a),
	.w7(32'h395629e9),
	.w8(32'h3b0818db),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a03d41e),
	.w1(32'hba2a7ffe),
	.w2(32'hb9471334),
	.w3(32'h39d9ce30),
	.w4(32'hb98b0489),
	.w5(32'h3a0188b5),
	.w6(32'hbaa16321),
	.w7(32'hba66b8dc),
	.w8(32'h39a09d90),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a906717),
	.w1(32'hb918e53a),
	.w2(32'h3a0382e7),
	.w3(32'h3a99d46b),
	.w4(32'h3ae29acb),
	.w5(32'h3ab78c1c),
	.w6(32'h3a1a8a46),
	.w7(32'h3a4fde7d),
	.w8(32'h3b1a6e62),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0d8a7c),
	.w1(32'h39d4cd0e),
	.w2(32'h3a4b013a),
	.w3(32'h3b5acc3e),
	.w4(32'hb9873cdb),
	.w5(32'hba58e351),
	.w6(32'h3ac29a5f),
	.w7(32'hb70f2f5c),
	.w8(32'hba81a92c),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaddf97d),
	.w1(32'h3b098a51),
	.w2(32'h37aac6d6),
	.w3(32'hbaa75bfb),
	.w4(32'h3acf9c7f),
	.w5(32'hba10668d),
	.w6(32'h3b04fc82),
	.w7(32'hba4444dd),
	.w8(32'hb9cb7322),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba66f0ab),
	.w1(32'h3abcb51e),
	.w2(32'h3b5124e8),
	.w3(32'hba814a65),
	.w4(32'hb9ac7774),
	.w5(32'hba859923),
	.w6(32'h3a98af23),
	.w7(32'h3b19a2c7),
	.w8(32'hb7f4dd32),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4c903c),
	.w1(32'hba97f24c),
	.w2(32'h3b26723d),
	.w3(32'hbb7abaf8),
	.w4(32'hba3b0e0b),
	.w5(32'h3b50503e),
	.w6(32'hbad3d10e),
	.w7(32'h3b206e32),
	.w8(32'h3b0f234e),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2e6e59),
	.w1(32'h39862ac7),
	.w2(32'h39b3624b),
	.w3(32'h39beb076),
	.w4(32'h3a327862),
	.w5(32'hb79ce32a),
	.w6(32'hb975a89f),
	.w7(32'hb8c941bf),
	.w8(32'hba9b6e75),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadecbc2),
	.w1(32'h3b7a5330),
	.w2(32'h3ab3ad65),
	.w3(32'hbacdbce4),
	.w4(32'h3b5fc503),
	.w5(32'h39a0187f),
	.w6(32'h3b60f008),
	.w7(32'h3a211a33),
	.w8(32'h3a151e6f),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ca3329),
	.w1(32'hbaa0c682),
	.w2(32'hbb249220),
	.w3(32'h38310520),
	.w4(32'hba8d8f39),
	.w5(32'hbabc4535),
	.w6(32'hbae58b94),
	.w7(32'hbb0a5bbb),
	.w8(32'hba2936d9),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba15f9c7),
	.w1(32'h3a1feeab),
	.w2(32'hb95ac68a),
	.w3(32'hba1b795c),
	.w4(32'hbaa5c336),
	.w5(32'hb9c45681),
	.w6(32'h3a19b432),
	.w7(32'hb83568a4),
	.w8(32'hba5502a6),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b834e6),
	.w1(32'h3ba6c734),
	.w2(32'h3a710fb3),
	.w3(32'hb9cc79e3),
	.w4(32'h3b198790),
	.w5(32'hba7c6731),
	.w6(32'h3b186b68),
	.w7(32'hbb055225),
	.w8(32'hbac88293),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7747b7),
	.w1(32'hb9c57de0),
	.w2(32'hbad058a1),
	.w3(32'hbb8bcca7),
	.w4(32'h39b30fab),
	.w5(32'hba786f06),
	.w6(32'h3a138860),
	.w7(32'hbaf0d8ee),
	.w8(32'hba6e9261),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c57688),
	.w1(32'h3aab14bd),
	.w2(32'h38eed2e0),
	.w3(32'h3a6a110a),
	.w4(32'h3ae1f898),
	.w5(32'h3a35a9ce),
	.w6(32'h3b3af359),
	.w7(32'hba7b8826),
	.w8(32'hb9739bb3),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89d3d1c),
	.w1(32'hbb499454),
	.w2(32'hba8a800f),
	.w3(32'h39ef183b),
	.w4(32'hbb20e6e2),
	.w5(32'hbb3a1d37),
	.w6(32'hbb44fbdf),
	.w7(32'hb6e9fa8c),
	.w8(32'h382db1c4),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3a40e2),
	.w1(32'h3b35b90a),
	.w2(32'h3a6079b3),
	.w3(32'hba014c7a),
	.w4(32'h3b14b80c),
	.w5(32'h399f237b),
	.w6(32'h3b13e4d3),
	.w7(32'h3800a4a5),
	.w8(32'h3a980327),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a585712),
	.w1(32'h39e18983),
	.w2(32'hbaa039df),
	.w3(32'h3a5abf5e),
	.w4(32'h3ace25b5),
	.w5(32'hba6ca0b8),
	.w6(32'hba819b9b),
	.w7(32'hbb1952fc),
	.w8(32'h3a9c370c),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab8b635),
	.w1(32'h3c8a1b16),
	.w2(32'h3b007338),
	.w3(32'h3a96f8c1),
	.w4(32'h3c82a781),
	.w5(32'h3a9570aa),
	.w6(32'h3c7bd276),
	.w7(32'h3a381e90),
	.w8(32'hbafc49ce),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2c6e66),
	.w1(32'h3b0ab896),
	.w2(32'h3a7aac1d),
	.w3(32'hbab500d9),
	.w4(32'h39d26466),
	.w5(32'h3942c92b),
	.w6(32'h3b8f3a7e),
	.w7(32'h3b836602),
	.w8(32'h3b905554),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af4b4eb),
	.w1(32'h3a4bb13a),
	.w2(32'hb97b493a),
	.w3(32'h38890e19),
	.w4(32'h3a9c8364),
	.w5(32'h3999ea76),
	.w6(32'h3a06ddf2),
	.w7(32'hb9cdcf58),
	.w8(32'hb8f462aa),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3822d156),
	.w1(32'h3a58b040),
	.w2(32'h38d8bb68),
	.w3(32'h38c89889),
	.w4(32'h3a8fde00),
	.w5(32'h388f988e),
	.w6(32'h3994e2e8),
	.w7(32'hba65fb52),
	.w8(32'h392f6ea3),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9fd2d0),
	.w1(32'h3aa8b803),
	.w2(32'h3a339242),
	.w3(32'h3a9f7825),
	.w4(32'h3ab18ca5),
	.w5(32'hb96457f2),
	.w6(32'h3919490b),
	.w7(32'hba82744b),
	.w8(32'h3a3b35c9),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a940ba9),
	.w1(32'h3bce8c35),
	.w2(32'h3bae13e9),
	.w3(32'h39dc8b1d),
	.w4(32'h3c17d02f),
	.w5(32'h3bf0ee5e),
	.w6(32'h3bf9c8cf),
	.w7(32'h3b8f72bc),
	.w8(32'h3b402b4b),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9e49a7),
	.w1(32'hba2c1701),
	.w2(32'h3a27e530),
	.w3(32'h3b5b8ccd),
	.w4(32'h392b59b4),
	.w5(32'h3aa3bfdb),
	.w6(32'hb98e1c7a),
	.w7(32'h3a6cf869),
	.w8(32'h3b1247cb),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af02059),
	.w1(32'h3a42c17e),
	.w2(32'h3955edda),
	.w3(32'h3b040364),
	.w4(32'h382ef480),
	.w5(32'hba7992c3),
	.w6(32'h39e33fd9),
	.w7(32'hba811376),
	.w8(32'h393a0896),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb95e621c),
	.w1(32'hbb230d7e),
	.w2(32'h3b297020),
	.w3(32'hb8dd4763),
	.w4(32'hbb0389f2),
	.w5(32'h3b2714f5),
	.w6(32'hbb018d4a),
	.w7(32'h39922f82),
	.w8(32'h3a1fe135),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8a1e32),
	.w1(32'hbaf3554d),
	.w2(32'hb84a3a1c),
	.w3(32'h39e2fa82),
	.w4(32'hbb157e8f),
	.w5(32'hba29bdf3),
	.w6(32'h3a7e40ec),
	.w7(32'h39671cf7),
	.w8(32'hba8539ba),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb84776be),
	.w1(32'h387bf5f2),
	.w2(32'hbaf5fb87),
	.w3(32'hb956a958),
	.w4(32'h39b6c04c),
	.w5(32'hbadcfe86),
	.w6(32'h3aad7ddb),
	.w7(32'hbb0901e6),
	.w8(32'hbadeaac6),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba62725d),
	.w1(32'hbb1737a9),
	.w2(32'hba82c3a2),
	.w3(32'hb9acbd52),
	.w4(32'hbb160824),
	.w5(32'hba878645),
	.w6(32'hbaba0a35),
	.w7(32'hba4a01f2),
	.w8(32'hbac715bd),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaa4d8c),
	.w1(32'h3b915b85),
	.w2(32'h3614e6ae),
	.w3(32'hbae254d0),
	.w4(32'h3b94d880),
	.w5(32'h3a2bc8a4),
	.w6(32'h3bb12066),
	.w7(32'h3b6705aa),
	.w8(32'h3b88954e),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab300ad),
	.w1(32'h38a0b8c2),
	.w2(32'h3abaf349),
	.w3(32'h3a022d74),
	.w4(32'hbae66b84),
	.w5(32'hba5365f8),
	.w6(32'hba4b7927),
	.w7(32'h3a1a4ec9),
	.w8(32'h38cee325),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9148e14),
	.w1(32'hba205f9f),
	.w2(32'hba0bd28a),
	.w3(32'hbae6c520),
	.w4(32'hb9aec68f),
	.w5(32'hba0d4e6b),
	.w6(32'hb9db81bd),
	.w7(32'hbabec91c),
	.w8(32'hb880402f),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4e3f5d),
	.w1(32'h3a2b2416),
	.w2(32'h3ab2d279),
	.w3(32'h3a52804a),
	.w4(32'h3b24f44d),
	.w5(32'h3b5d8b6e),
	.w6(32'h3b31d0a9),
	.w7(32'h3ba9cdf9),
	.w8(32'h3ba19764),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa24403),
	.w1(32'hbac89729),
	.w2(32'h39b5026c),
	.w3(32'h3b4625ee),
	.w4(32'hb9cc8cb6),
	.w5(32'h39dd85bb),
	.w6(32'hb999a057),
	.w7(32'h3a9b5e1b),
	.w8(32'h3a37e164),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38bee6b1),
	.w1(32'hba5df066),
	.w2(32'hb968d843),
	.w3(32'hb9a80fd1),
	.w4(32'hba0ce57f),
	.w5(32'h3947efb4),
	.w6(32'h38e17efd),
	.w7(32'hb9dd46f0),
	.w8(32'h3a046a89),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa42982),
	.w1(32'h3aaadd65),
	.w2(32'hb96c5f1d),
	.w3(32'h3ac2991b),
	.w4(32'h3af53dda),
	.w5(32'h3b1f622d),
	.w6(32'h3acba0b9),
	.w7(32'h3a239fdd),
	.w8(32'hba39f0ad),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb51a4d1),
	.w1(32'h3cb41f80),
	.w2(32'h3c3d0501),
	.w3(32'hba028e4c),
	.w4(32'h3c956882),
	.w5(32'h3c0a4ea6),
	.w6(32'h3c8c68b9),
	.w7(32'h3bfdaaa7),
	.w8(32'h3ae9724e),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b526e1c),
	.w1(32'hb9838b69),
	.w2(32'h386eb117),
	.w3(32'hbab48000),
	.w4(32'h3908a9ee),
	.w5(32'hb9d08e94),
	.w6(32'hb9a212f4),
	.w7(32'hba9e8b66),
	.w8(32'h39ae4943),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa465cb),
	.w1(32'h37f19331),
	.w2(32'hba54b53f),
	.w3(32'h3a467ea1),
	.w4(32'h3a572f02),
	.w5(32'h38bde88f),
	.w6(32'h39a729a3),
	.w7(32'hba22ddc0),
	.w8(32'hb9d1ca8e),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d5e9e2),
	.w1(32'h3aefb03d),
	.w2(32'h3a90c6ef),
	.w3(32'h3a0acc91),
	.w4(32'h3acace6c),
	.w5(32'h3a93ddd4),
	.w6(32'h3a9ee462),
	.w7(32'h3a490dd6),
	.w8(32'hb9956bf2),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb638c5d8),
	.w1(32'h3baa3678),
	.w2(32'hba9ad80c),
	.w3(32'h3a8c6228),
	.w4(32'h3b8e7972),
	.w5(32'hbacff132),
	.w6(32'h3b5ba935),
	.w7(32'hba78c857),
	.w8(32'h3af0b986),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a02d9a5),
	.w1(32'h3aa106e5),
	.w2(32'h3a20f343),
	.w3(32'h3b0858c4),
	.w4(32'h39c76fbc),
	.w5(32'hba864a99),
	.w6(32'h3abd84d1),
	.w7(32'hb9f16284),
	.w8(32'h3ada1c56),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6c5eee),
	.w1(32'hba7023ff),
	.w2(32'h39a273f2),
	.w3(32'hba1f1558),
	.w4(32'h398a5d41),
	.w5(32'h3a2d08ab),
	.w6(32'hb9d06943),
	.w7(32'h3a9763a4),
	.w8(32'hba4a8214),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba623ecb),
	.w1(32'hba08c0fb),
	.w2(32'hba28abff),
	.w3(32'hba8a0139),
	.w4(32'hba026088),
	.w5(32'hb9f250ee),
	.w6(32'hb9b66641),
	.w7(32'hb9c48d36),
	.w8(32'hb8562afd),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dbd1e7),
	.w1(32'h3959b206),
	.w2(32'h38fc8c03),
	.w3(32'hba1874fe),
	.w4(32'h3a82a822),
	.w5(32'h3a4b219a),
	.w6(32'h3ad71392),
	.w7(32'h3b219139),
	.w8(32'h3b8ecf64),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af064de),
	.w1(32'h39e33fbb),
	.w2(32'hb92266d4),
	.w3(32'h3af520eb),
	.w4(32'h3a6decde),
	.w5(32'hb990f344),
	.w6(32'h3a46011c),
	.w7(32'h396b4ce6),
	.w8(32'hb9d1266e),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0e9d68),
	.w1(32'h3a79cc48),
	.w2(32'hbb19b36b),
	.w3(32'hbab56bc7),
	.w4(32'h3a3b618a),
	.w5(32'hbb0182bc),
	.w6(32'h3a95d309),
	.w7(32'hbad151f6),
	.w8(32'hba899cd0),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1cf3db),
	.w1(32'hb9c1ec62),
	.w2(32'hba5132b8),
	.w3(32'h3a0549c5),
	.w4(32'hb8ea6819),
	.w5(32'hba0b85f2),
	.w6(32'hb6b16d98),
	.w7(32'hba0c082a),
	.w8(32'hbad1b8af),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabbcc63),
	.w1(32'h398af564),
	.w2(32'hbad897f7),
	.w3(32'hba8ad564),
	.w4(32'h3a65d219),
	.w5(32'hba96b445),
	.w6(32'h39a3937d),
	.w7(32'hbb002ece),
	.w8(32'hba864ae1),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba82cafe),
	.w1(32'hbb0004ec),
	.w2(32'hbab2849b),
	.w3(32'hb99c4aac),
	.w4(32'hbb083168),
	.w5(32'hbace43c3),
	.w6(32'hbb0dc6c4),
	.w7(32'hbaa6824c),
	.w8(32'hbaa1e458),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad21772),
	.w1(32'h374bf893),
	.w2(32'hba4c1b43),
	.w3(32'hbb17aec3),
	.w4(32'h3a89a00b),
	.w5(32'hb795355d),
	.w6(32'hba3747bd),
	.w7(32'hba209803),
	.w8(32'h3a35461e),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fabdbe),
	.w1(32'h3bd30f09),
	.w2(32'h3b708fa7),
	.w3(32'hb71321de),
	.w4(32'h3bbdaa10),
	.w5(32'h3b31d661),
	.w6(32'h3b84ef38),
	.w7(32'h3ac40872),
	.w8(32'h3b317aac),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1c224c),
	.w1(32'h387b4282),
	.w2(32'h3a21bb6d),
	.w3(32'hb9d5d4f9),
	.w4(32'h3a842e0d),
	.w5(32'h3ae98182),
	.w6(32'h3acb49dc),
	.w7(32'h3b39d3f2),
	.w8(32'h3b31c945),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a404d1d),
	.w1(32'hbb0abefa),
	.w2(32'hbadf8b1f),
	.w3(32'h3ad34618),
	.w4(32'hba9fc4c5),
	.w5(32'hba4d00c1),
	.w6(32'hbabe90f3),
	.w7(32'hbac57dc8),
	.w8(32'hb9426e17),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a017cc4),
	.w1(32'h39c29f40),
	.w2(32'hba99dc8e),
	.w3(32'h38ee6f7a),
	.w4(32'h3a1a7e91),
	.w5(32'hba0036aa),
	.w6(32'h3a4979e5),
	.w7(32'hb8959abf),
	.w8(32'hb9e3e82f),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a828e3a),
	.w1(32'h3bc88755),
	.w2(32'h3be15b3b),
	.w3(32'h3aab397f),
	.w4(32'h3bd185e6),
	.w5(32'h3b9a9d0d),
	.w6(32'h3be2bde4),
	.w7(32'h3c03577b),
	.w8(32'h3c163ebf),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc519ef),
	.w1(32'h3bd5325f),
	.w2(32'hbafc805f),
	.w3(32'h3b9a4f6f),
	.w4(32'h3be509e2),
	.w5(32'hb851e724),
	.w6(32'h3c04f308),
	.w7(32'h3a181ed3),
	.w8(32'h39b94672),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb979ea2b),
	.w1(32'h3a09c298),
	.w2(32'hba09570a),
	.w3(32'hbb281446),
	.w4(32'h39fb3af3),
	.w5(32'hba41c29d),
	.w6(32'h3988f4cc),
	.w7(32'hba863d53),
	.w8(32'h37021d24),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba700afe),
	.w1(32'hba4bef28),
	.w2(32'hb8c6f7d3),
	.w3(32'hb9a91aa6),
	.w4(32'h391ee945),
	.w5(32'h3b20db7a),
	.w6(32'h3aa41835),
	.w7(32'h398bf8ed),
	.w8(32'hb92e1876),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa111d9),
	.w1(32'hba5290e0),
	.w2(32'h3ab1a46f),
	.w3(32'h3b6f0786),
	.w4(32'hba189ea1),
	.w5(32'h3a4d021e),
	.w6(32'hba11a26b),
	.w7(32'h3aad34f0),
	.w8(32'h39cdd897),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3979ac07),
	.w1(32'hb930c6d4),
	.w2(32'hbab0be4e),
	.w3(32'hb8f2969a),
	.w4(32'h3985a506),
	.w5(32'hba4fd0fe),
	.w6(32'h375bb00e),
	.w7(32'hbac6be0b),
	.w8(32'hba410fb8),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0326f3),
	.w1(32'h39aee4f8),
	.w2(32'hbacd35ea),
	.w3(32'hb7ee0ffa),
	.w4(32'h3a2f850f),
	.w5(32'hba9b96fd),
	.w6(32'h39ba1aa3),
	.w7(32'hbae70d4e),
	.w8(32'hba7b2986),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba88a3b3),
	.w1(32'h3a885458),
	.w2(32'h37c1467c),
	.w3(32'hba0e88cb),
	.w4(32'h3a86f40a),
	.w5(32'hb9572fb4),
	.w6(32'h395b8ddd),
	.w7(32'hbac765b2),
	.w8(32'hb8f98f4e),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abce6fe),
	.w1(32'h3a13e81d),
	.w2(32'hb77bcb51),
	.w3(32'h3a832e51),
	.w4(32'h39c876e5),
	.w5(32'hba72d111),
	.w6(32'h39ce3d25),
	.w7(32'hb997afcc),
	.w8(32'hba87265a),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad50e3b),
	.w1(32'hbad195be),
	.w2(32'h3a99f88c),
	.w3(32'hbac908f5),
	.w4(32'hbb908d14),
	.w5(32'hbb4021ac),
	.w6(32'hbb6cb24c),
	.w7(32'h3a955a00),
	.w8(32'h3b104434),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf872dd),
	.w1(32'h3a965f2f),
	.w2(32'hba12965f),
	.w3(32'hbafb3fdc),
	.w4(32'h3b3b1773),
	.w5(32'h3ab040ce),
	.w6(32'h3b1850db),
	.w7(32'hb92b3f19),
	.w8(32'h3b13ecd8),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae49a36),
	.w1(32'h3b41e1f0),
	.w2(32'h3ad37344),
	.w3(32'h3b4b911f),
	.w4(32'h3b50be01),
	.w5(32'h3a43d300),
	.w6(32'h3b246f4d),
	.w7(32'h3aa9d89a),
	.w8(32'hba7213b0),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabb1383),
	.w1(32'hbb1f9d4e),
	.w2(32'hba29f905),
	.w3(32'hbad1a051),
	.w4(32'hbb534c77),
	.w5(32'hbb66ef87),
	.w6(32'hbb05b782),
	.w7(32'hb98b52d6),
	.w8(32'hba0442f8),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba959548),
	.w1(32'h3b1e0091),
	.w2(32'hba083e59),
	.w3(32'hbb02fb67),
	.w4(32'h3b3303a2),
	.w5(32'h3914aac1),
	.w6(32'h3b0b94cb),
	.w7(32'hba14e7df),
	.w8(32'hb9d26ac9),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb982b0b2),
	.w1(32'h3c3a0d5f),
	.w2(32'h3b80a1a5),
	.w3(32'h38a842d1),
	.w4(32'h3c34f39b),
	.w5(32'h3b82fb6f),
	.w6(32'h3c3fabea),
	.w7(32'h3b9f5af9),
	.w8(32'h3b482b4b),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b24031f),
	.w1(32'hba640513),
	.w2(32'h3ae28c08),
	.w3(32'hb99a2efb),
	.w4(32'hbaa9b1c2),
	.w5(32'h3a9a8154),
	.w6(32'hba88f75c),
	.w7(32'h3a99fbc7),
	.w8(32'h39b26bf0),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37009129),
	.w1(32'h3ba447b1),
	.w2(32'h3b2895bd),
	.w3(32'hba5f6d4b),
	.w4(32'h3b4fb264),
	.w5(32'h38ae9480),
	.w6(32'h3b8d4fa7),
	.w7(32'h3aedbce7),
	.w8(32'h3a84c803),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a13690f),
	.w1(32'hba861f7d),
	.w2(32'hb978e36f),
	.w3(32'hba15aa3e),
	.w4(32'hbacd0c90),
	.w5(32'hba2a2c2c),
	.w6(32'hba300bb5),
	.w7(32'hb9a5d8ae),
	.w8(32'hbac8f05f),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab19f4a),
	.w1(32'h3c251a14),
	.w2(32'h3c3433c5),
	.w3(32'hbad7698d),
	.w4(32'h3bbb18e3),
	.w5(32'h3bc7cc77),
	.w6(32'h3bd35588),
	.w7(32'h3b32f70a),
	.w8(32'hb96b0d7e),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfc4b07),
	.w1(32'h3ad3719e),
	.w2(32'h3ba55918),
	.w3(32'hbabcfd7a),
	.w4(32'h3a76b5f6),
	.w5(32'h3b5f5dab),
	.w6(32'h3b00abd8),
	.w7(32'h3ba6b347),
	.w8(32'h3b20e1bd),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1305fd),
	.w1(32'hb90d056f),
	.w2(32'h3b24d9b0),
	.w3(32'h3a7da7d5),
	.w4(32'h3a803b55),
	.w5(32'h3b02fffa),
	.w6(32'hb879e638),
	.w7(32'h3ab8c2f6),
	.w8(32'h3aa231f0),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2bad9a),
	.w1(32'h39b4f8e3),
	.w2(32'hba594f2e),
	.w3(32'h3b2d0e2f),
	.w4(32'h3a1e3e8e),
	.w5(32'hb981b905),
	.w6(32'h3915a42e),
	.w7(32'hba809b65),
	.w8(32'hb99f716b),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88ea78e),
	.w1(32'hb8e30ed5),
	.w2(32'hba57622b),
	.w3(32'h39c3e0a5),
	.w4(32'hb87f2d52),
	.w5(32'hba0d4320),
	.w6(32'h3a6af849),
	.w7(32'hb92fc312),
	.w8(32'h39989cfe),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba395421),
	.w1(32'h3a53e18e),
	.w2(32'hba358be0),
	.w3(32'hb9fea7d3),
	.w4(32'h3aeea806),
	.w5(32'h3a314a22),
	.w6(32'h3a479503),
	.w7(32'hba07e280),
	.w8(32'h3a93338e),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3991ee59),
	.w1(32'hb9a13efc),
	.w2(32'hba0645af),
	.w3(32'h3a53a760),
	.w4(32'h39b9f579),
	.w5(32'hb9460e9b),
	.w6(32'hba6c1895),
	.w7(32'hbb03d81e),
	.w8(32'hba290390),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39296116),
	.w1(32'hb9c6483c),
	.w2(32'h3b0c34dd),
	.w3(32'h39decf32),
	.w4(32'hba27d1a5),
	.w5(32'h3aa591bb),
	.w6(32'h39c10548),
	.w7(32'h3b2fadb8),
	.w8(32'h3ae88d8a),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39aa1c9d),
	.w1(32'hba6905a3),
	.w2(32'h3afb9cb2),
	.w3(32'hb9dbda63),
	.w4(32'hbae901c6),
	.w5(32'h3a1abada),
	.w6(32'h37c21dcb),
	.w7(32'h3ab3100d),
	.w8(32'h3b0c2860),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0d0be6),
	.w1(32'h3bd182f9),
	.w2(32'hbac0da05),
	.w3(32'h39c88333),
	.w4(32'h3bce2f91),
	.w5(32'h388ab808),
	.w6(32'h3bda8047),
	.w7(32'h3841e247),
	.w8(32'h35a9fb65),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b89ff9),
	.w1(32'hba55ed95),
	.w2(32'h37a47adb),
	.w3(32'hba8c9547),
	.w4(32'hbac26f83),
	.w5(32'hba564547),
	.w6(32'hba632b61),
	.w7(32'hbaa419a8),
	.w8(32'hbaefe6a0),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba20447f),
	.w1(32'hbaa2dbc4),
	.w2(32'h399a01af),
	.w3(32'hbab50449),
	.w4(32'hbacf3a01),
	.w5(32'h3aaba96d),
	.w6(32'hb811fe2f),
	.w7(32'hb9277fb0),
	.w8(32'hba0dda9d),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad8e82c),
	.w1(32'h3bf8260c),
	.w2(32'h3abe6065),
	.w3(32'h3b0cb4c3),
	.w4(32'h3bc2f558),
	.w5(32'h3a4bd5e2),
	.w6(32'h3bbc842a),
	.w7(32'h39eed947),
	.w8(32'hbb1a96e3),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae16cb8),
	.w1(32'h3b30fc6f),
	.w2(32'hbb1f05e8),
	.w3(32'hbba4dade),
	.w4(32'h3b9f7b8e),
	.w5(32'hbaaa2c5a),
	.w6(32'h3b3ea7b7),
	.w7(32'hbada1dec),
	.w8(32'h3b4c6b43),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2f4bb4),
	.w1(32'hbaecf022),
	.w2(32'h3a54d2e7),
	.w3(32'h3ae64d3b),
	.w4(32'hbb1070da),
	.w5(32'h3a28e7f6),
	.w6(32'hbb0167d5),
	.w7(32'h3857de89),
	.w8(32'hba8bc40f),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabd4218),
	.w1(32'h3b2f2b77),
	.w2(32'h3b3a791d),
	.w3(32'hba89a688),
	.w4(32'h3b1712e7),
	.w5(32'h3b06e1d8),
	.w6(32'h3b81ae8b),
	.w7(32'h3a953016),
	.w8(32'h3b73afbc),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1e2032),
	.w1(32'h3aaca6b1),
	.w2(32'hbb1137bf),
	.w3(32'h3a718829),
	.w4(32'h3a93c9e6),
	.w5(32'hbb1da557),
	.w6(32'h3b8dda78),
	.w7(32'hbb18cb78),
	.w8(32'hbad52a60),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0c7e78),
	.w1(32'hb94f671e),
	.w2(32'hba05576b),
	.w3(32'h3b142f4d),
	.w4(32'hbac588d9),
	.w5(32'hbaf1b76c),
	.w6(32'h3a4f03ea),
	.w7(32'h3a91c0a6),
	.w8(32'hba994e96),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaafb3ce),
	.w1(32'h3ac4e813),
	.w2(32'hba871c9f),
	.w3(32'hbaa54284),
	.w4(32'h3b6e7420),
	.w5(32'h3aca2e48),
	.w6(32'h3b2a01fa),
	.w7(32'hba414cc0),
	.w8(32'h3b48c6b4),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b163836),
	.w1(32'h38a106bd),
	.w2(32'hbaa98feb),
	.w3(32'h3b889908),
	.w4(32'h3a0d6175),
	.w5(32'hba3b8377),
	.w6(32'h39808ab3),
	.w7(32'hbaa32f2a),
	.w8(32'hb9d3780c),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b09cdf),
	.w1(32'h3a43b569),
	.w2(32'h3a093299),
	.w3(32'h38897c30),
	.w4(32'h3b16602b),
	.w5(32'h3b003e8f),
	.w6(32'h3b0f5149),
	.w7(32'hb9bdff75),
	.w8(32'h3b134b8c),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1f2311),
	.w1(32'h3b1a78fe),
	.w2(32'h3ac89eb6),
	.w3(32'h3ae839a9),
	.w4(32'h3b0c6f32),
	.w5(32'h39e7c455),
	.w6(32'h3b1a6de7),
	.w7(32'h39d2a08e),
	.w8(32'h3a7b87d2),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a456c2a),
	.w1(32'hba7e4b16),
	.w2(32'hba88189c),
	.w3(32'h3a08e94b),
	.w4(32'hbb210b04),
	.w5(32'hbb0385b5),
	.w6(32'hbacd4976),
	.w7(32'hbb176155),
	.w8(32'hbb2f7945),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad154b6),
	.w1(32'hba0d0af3),
	.w2(32'hbab1a00d),
	.w3(32'hbb30810e),
	.w4(32'hb9b71765),
	.w5(32'hba161f38),
	.w6(32'hbadef8c6),
	.w7(32'hbb168a91),
	.w8(32'hba9a837b),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98370b5),
	.w1(32'h3a446c86),
	.w2(32'hba331cc4),
	.w3(32'hb9a901ad),
	.w4(32'h3afeb36f),
	.w5(32'h3a33099b),
	.w6(32'h3ac53a7b),
	.w7(32'hb6ae5054),
	.w8(32'h3ad22233),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab7bda6),
	.w1(32'hbb7f721c),
	.w2(32'hbb09b3af),
	.w3(32'h3b2de1d1),
	.w4(32'hbb554e59),
	.w5(32'hbb1f129f),
	.w6(32'hbb4e8897),
	.w7(32'hbb3a33c3),
	.w8(32'hbb3faa03),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2e3cef),
	.w1(32'h3ac31391),
	.w2(32'hba633370),
	.w3(32'hbb611499),
	.w4(32'h3aaed676),
	.w5(32'hbac55f58),
	.w6(32'h3ae1bd73),
	.w7(32'hbaab8eaa),
	.w8(32'hb9af6ecb),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cd1ddf),
	.w1(32'h3ab68fb1),
	.w2(32'hb8262b79),
	.w3(32'hb91cd8bd),
	.w4(32'h3b23bb44),
	.w5(32'hba6fd24b),
	.w6(32'h3aac75a2),
	.w7(32'hba00770c),
	.w8(32'h3b545890),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8a622c),
	.w1(32'h3b38d96d),
	.w2(32'h390be856),
	.w3(32'h3a6cfa60),
	.w4(32'h3b125e49),
	.w5(32'hba69fdc9),
	.w6(32'h3b560850),
	.w7(32'hba304e98),
	.w8(32'h39836b55),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94edc20),
	.w1(32'hbaad8c15),
	.w2(32'hba94c685),
	.w3(32'hb9f6bfc9),
	.w4(32'hbacc0222),
	.w5(32'hbafede49),
	.w6(32'hbb112b90),
	.w7(32'hbaf85003),
	.w8(32'hbb045b66),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0368d3),
	.w1(32'hbb41c4e7),
	.w2(32'hbabd5f9a),
	.w3(32'hbb03e19d),
	.w4(32'hbae1268b),
	.w5(32'hbad65d78),
	.w6(32'hbabd101a),
	.w7(32'hbaf1180a),
	.w8(32'h3903243b),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3954133e),
	.w1(32'h3aaba82d),
	.w2(32'hba86e63e),
	.w3(32'hba6506a0),
	.w4(32'h3b36d02e),
	.w5(32'h3a2820f8),
	.w6(32'h3b1a6b9a),
	.w7(32'hb89813f3),
	.w8(32'h3b048312),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae8252c),
	.w1(32'hb9f76356),
	.w2(32'hba947aec),
	.w3(32'h3b4d5ce8),
	.w4(32'hb98498c0),
	.w5(32'hba5c5fdb),
	.w6(32'h377b1e77),
	.w7(32'hba67b696),
	.w8(32'h3935dedb),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396d5cd0),
	.w1(32'hb8851e74),
	.w2(32'hbaad1758),
	.w3(32'h399319af),
	.w4(32'h3900e3f1),
	.w5(32'hba7fdd2a),
	.w6(32'h3a050000),
	.w7(32'hba8b222b),
	.w8(32'h39839137),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a79fae),
	.w1(32'hbaa3066c),
	.w2(32'hba9a4aeb),
	.w3(32'h3a1878f6),
	.w4(32'hba81d6b4),
	.w5(32'hb9c64615),
	.w6(32'hbaad81d1),
	.w7(32'hbad364b4),
	.w8(32'h38e7fd77),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a040daa),
	.w1(32'h3b4101e8),
	.w2(32'hbaeb3ab4),
	.w3(32'h3a0dd767),
	.w4(32'h3b4e4b52),
	.w5(32'hbad38eb9),
	.w6(32'h3b7c43a7),
	.w7(32'hba8bd7f8),
	.w8(32'hbb2b875e),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb032ca1),
	.w1(32'h3b0159e9),
	.w2(32'h3a2259fb),
	.w3(32'hbb12b94a),
	.w4(32'h3aecf987),
	.w5(32'h37e259fd),
	.w6(32'h3b01779b),
	.w7(32'hba2cdd90),
	.w8(32'h3982b4a4),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4898c5),
	.w1(32'h3b548920),
	.w2(32'h3a7cd154),
	.w3(32'hb9a1318c),
	.w4(32'h3b3aaf50),
	.w5(32'h39acb862),
	.w6(32'h3b11894a),
	.w7(32'hb9de8da2),
	.w8(32'hb9b07305),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba15f404),
	.w1(32'hba045824),
	.w2(32'hbaf22aa1),
	.w3(32'hba2158fa),
	.w4(32'h390d745e),
	.w5(32'hba9e5c80),
	.w6(32'h3a835a22),
	.w7(32'hbafb0c65),
	.w8(32'hba6dce96),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba56ed85),
	.w1(32'h3aaca624),
	.w2(32'hbacd7ab8),
	.w3(32'h383bd40e),
	.w4(32'hba778c21),
	.w5(32'hbb4e51aa),
	.w6(32'h3ab3bae9),
	.w7(32'h399ce54e),
	.w8(32'hb9f3f579),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba93634c),
	.w1(32'h3a93cbcb),
	.w2(32'h3ab28104),
	.w3(32'hbafa53c5),
	.w4(32'hb9225e56),
	.w5(32'h38e68c03),
	.w6(32'h3afd3440),
	.w7(32'h39d933a4),
	.w8(32'h3ae2bf5f),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2309ca),
	.w1(32'h3b91341b),
	.w2(32'hb99eacf1),
	.w3(32'h379accba),
	.w4(32'h3b84e676),
	.w5(32'hb94d379f),
	.w6(32'h3b6e759f),
	.w7(32'hba4dc9eb),
	.w8(32'hb80f00d1),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c9d8cd),
	.w1(32'hb87ba9b0),
	.w2(32'hb8658564),
	.w3(32'h3989d3be),
	.w4(32'hb8dfbd39),
	.w5(32'hb8ca3aac),
	.w6(32'hb8209d1d),
	.w7(32'hb83e8f95),
	.w8(32'hb88b070f),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba05f0a0),
	.w1(32'hb817e7d6),
	.w2(32'h38679c6e),
	.w3(32'hb9cb19b7),
	.w4(32'h38c7e1b6),
	.w5(32'h3915fc16),
	.w6(32'h38105fb6),
	.w7(32'h38808db5),
	.w8(32'h3a001a2a),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96322c8),
	.w1(32'h381ba335),
	.w2(32'h383066e8),
	.w3(32'hb7997ad9),
	.w4(32'h396fd4f5),
	.w5(32'h3927bf4a),
	.w6(32'hb9569350),
	.w7(32'h38dcc5da),
	.w8(32'h39887e32),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb895afe5),
	.w1(32'hb5cbd5c4),
	.w2(32'h3838fa90),
	.w3(32'hb8006434),
	.w4(32'h3836c6d9),
	.w5(32'h38a3d24f),
	.w6(32'hb80bff40),
	.w7(32'hb6599d15),
	.w8(32'h38d74f02),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35dde529),
	.w1(32'hb8efef93),
	.w2(32'h37eaa84e),
	.w3(32'h38589e00),
	.w4(32'h36b5c3f6),
	.w5(32'h3891123b),
	.w6(32'h38e2a726),
	.w7(32'hb78ef9a0),
	.w8(32'h3877757d),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3744307b),
	.w1(32'hb89a4bd7),
	.w2(32'h38cd3708),
	.w3(32'h38bc23c1),
	.w4(32'hb80b0add),
	.w5(32'h38b00be0),
	.w6(32'h38df2780),
	.w7(32'hb719eeea),
	.w8(32'h38eff74f),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7369753),
	.w1(32'hb853cd99),
	.w2(32'hb7c40622),
	.w3(32'h3801bdc4),
	.w4(32'hb72c42de),
	.w5(32'h37c510c2),
	.w6(32'h383aa5db),
	.w7(32'h37d3b538),
	.w8(32'h38dbe03c),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3980e8fd),
	.w1(32'hb8594a22),
	.w2(32'h39b8bdd7),
	.w3(32'h395b4586),
	.w4(32'hb82faaa1),
	.w5(32'h38a9dabc),
	.w6(32'h39c1d85b),
	.w7(32'h3926d4d3),
	.w8(32'h394cd3ef),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba25f88c),
	.w1(32'h39a4f66f),
	.w2(32'h398ec999),
	.w3(32'hb91cef9c),
	.w4(32'h3a0d5df7),
	.w5(32'h3a1cf709),
	.w6(32'hb9637d1d),
	.w7(32'h396f43b2),
	.w8(32'h3a4627c3),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39063b48),
	.w1(32'hb9e882da),
	.w2(32'hb911c6ba),
	.w3(32'h39cd2d07),
	.w4(32'hb9b27407),
	.w5(32'hb90d4baf),
	.w6(32'h39cf9405),
	.w7(32'hb9530829),
	.w8(32'hb948a70d),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97cb306),
	.w1(32'hb8fc237b),
	.w2(32'h392ec315),
	.w3(32'hb9217b9a),
	.w4(32'hb91ed452),
	.w5(32'h39583fae),
	.w6(32'hb93a663c),
	.w7(32'hb940cc34),
	.w8(32'h395711f9),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d9c06a),
	.w1(32'h38ad62db),
	.w2(32'h392a89e2),
	.w3(32'hb930bd48),
	.w4(32'h39aeb790),
	.w5(32'h3a18de56),
	.w6(32'hb9062036),
	.w7(32'h3887ca08),
	.w8(32'h3a330be7),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d58b02),
	.w1(32'hba03b953),
	.w2(32'hb8159194),
	.w3(32'h37d606b0),
	.w4(32'hb9b731e2),
	.w5(32'hb799149c),
	.w6(32'h39a76600),
	.w7(32'hb8d29410),
	.w8(32'hb78fd6f6),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb958c4a3),
	.w1(32'hb8b160d5),
	.w2(32'h3701d8b8),
	.w3(32'h37aadd15),
	.w4(32'hb6881a70),
	.w5(32'h38d95483),
	.w6(32'hb8c05d21),
	.w7(32'hb8d30305),
	.w8(32'hb55f08da),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37e66ea0),
	.w1(32'hb7c846c0),
	.w2(32'h3812dd0a),
	.w3(32'h385c9457),
	.w4(32'h35fdaa83),
	.w5(32'h385d365c),
	.w6(32'h38780760),
	.w7(32'h380b81a7),
	.w8(32'h38e5b598),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a30e5b),
	.w1(32'hba7dce47),
	.w2(32'hba61e998),
	.w3(32'h3a1a0387),
	.w4(32'hb9b1a1ae),
	.w5(32'hba18966e),
	.w6(32'h3a1ff580),
	.w7(32'hb9ff72a1),
	.w8(32'hba0d3874),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb686db55),
	.w1(32'hb8f643fe),
	.w2(32'h39145b97),
	.w3(32'h38e3972f),
	.w4(32'h35df490f),
	.w5(32'h39827c01),
	.w6(32'h38f62a2a),
	.w7(32'hb854b14d),
	.w8(32'h3951bac4),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37203d26),
	.w1(32'h371e7e46),
	.w2(32'h370f8115),
	.w3(32'h371c5359),
	.w4(32'h372982d4),
	.w5(32'h37012363),
	.w6(32'hb4ed53ce),
	.w7(32'h368f930a),
	.w8(32'h351457b6),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5c94c10),
	.w1(32'hb719b771),
	.w2(32'hb64bd0e0),
	.w3(32'hb52619e2),
	.w4(32'hb68e2f09),
	.w5(32'hb6b963d4),
	.w6(32'h3736d3b7),
	.w7(32'h360d279a),
	.w8(32'h370ca789),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89c484f),
	.w1(32'hb93ffadc),
	.w2(32'h36f86f3a),
	.w3(32'hb7f289e1),
	.w4(32'hb90ccfc9),
	.w5(32'hb7d46f45),
	.w6(32'h38c4da79),
	.w7(32'hb8cf3f4d),
	.w8(32'hb806cea0),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h385c0f1e),
	.w1(32'hba301932),
	.w2(32'hb7c71fb8),
	.w3(32'h393c80cd),
	.w4(32'hba009950),
	.w5(32'h3892a777),
	.w6(32'h39ad5259),
	.w7(32'hb9f2f1fc),
	.w8(32'hb98e675f),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb881c3da),
	.w1(32'hb907f00b),
	.w2(32'h37fa70b6),
	.w3(32'h38b8c963),
	.w4(32'hb72a6c93),
	.w5(32'h3908697d),
	.w6(32'h38379d7b),
	.w7(32'h3816301e),
	.w8(32'h39fd5733),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb3ed0426),
	.w1(32'h33e9e1fa),
	.w2(32'hb54b69c5),
	.w3(32'hb4cab57c),
	.w4(32'hb554d503),
	.w5(32'hb655e43f),
	.w6(32'h355da71b),
	.w7(32'h358420e8),
	.w8(32'hb62a2ac2),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ad1de6),
	.w1(32'hb7b52b64),
	.w2(32'h38175126),
	.w3(32'h38f7802d),
	.w4(32'h3927771d),
	.w5(32'h3918921c),
	.w6(32'hb8a81b17),
	.w7(32'h381ce83d),
	.w8(32'h3950604a),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3798a950),
	.w1(32'hb968025b),
	.w2(32'hb87dc54a),
	.w3(32'h39262c21),
	.w4(32'hb8e1e061),
	.w5(32'h38255fbd),
	.w6(32'h38cdbd56),
	.w7(32'hb834f71f),
	.w8(32'h38350ee9),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b8705f),
	.w1(32'h394b75c5),
	.w2(32'h3986fe15),
	.w3(32'hb99b76c5),
	.w4(32'h38c80e17),
	.w5(32'h39ef92dd),
	.w6(32'hb9ea9ac5),
	.w7(32'hb9811b41),
	.w8(32'h39dabed4),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8250ca0),
	.w1(32'hb80ea84f),
	.w2(32'h38dd7d8c),
	.w3(32'h3997b341),
	.w4(32'h39498cf7),
	.w5(32'h390de0ed),
	.w6(32'h39c2bac8),
	.w7(32'h38f0bc96),
	.w8(32'h3863638f),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3883315e),
	.w1(32'hb91d362c),
	.w2(32'h38ba61d9),
	.w3(32'h38b75609),
	.w4(32'hb96e7bc8),
	.w5(32'hb7b8b47a),
	.w6(32'h38dd21a6),
	.w7(32'hb918f97c),
	.w8(32'hb814896f),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb86331fd),
	.w1(32'hb8bdcb19),
	.w2(32'hb7eea135),
	.w3(32'hb7d3d884),
	.w4(32'hb8a7e550),
	.w5(32'hb7a7b91f),
	.w6(32'hb6eac95c),
	.w7(32'hb8a2559a),
	.w8(32'hb7fbff96),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38f2f755),
	.w1(32'hb9b9cc99),
	.w2(32'hb8c7c32e),
	.w3(32'h3987d5c0),
	.w4(32'hb96cfadd),
	.w5(32'h37805441),
	.w6(32'h3992ad1d),
	.w7(32'hb92dc4ee),
	.w8(32'hb90173f9),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb883b5db),
	.w1(32'hb9df9fd8),
	.w2(32'h38836230),
	.w3(32'hb8865a1a),
	.w4(32'hba17cc3a),
	.w5(32'hb91308ae),
	.w6(32'hb86680ed),
	.w7(32'hb9feab26),
	.w8(32'hb8d676ad),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3928aaa1),
	.w1(32'hb94468df),
	.w2(32'h38327b19),
	.w3(32'h3914cc3d),
	.w4(32'hb97cffe4),
	.w5(32'hb814dad5),
	.w6(32'h39899a7e),
	.w7(32'hb90ddfaf),
	.w8(32'hb834d007),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a2caf4),
	.w1(32'h38081f36),
	.w2(32'h3890b321),
	.w3(32'h3878b00d),
	.w4(32'h392760d4),
	.w5(32'h393dfe04),
	.w6(32'hb80eb45d),
	.w7(32'h36b85a34),
	.w8(32'h395e42a7),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37a67ccf),
	.w1(32'h352f9c38),
	.w2(32'h37ae6241),
	.w3(32'h381fe5a1),
	.w4(32'hb611529b),
	.w5(32'h37b49497),
	.w6(32'h378ca7be),
	.w7(32'h35c5ea38),
	.w8(32'hb6f1a2b3),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94d695f),
	.w1(32'hb84df899),
	.w2(32'h33fd7b18),
	.w3(32'h38232ef9),
	.w4(32'h386b9a36),
	.w5(32'h3918ef4f),
	.w6(32'h38100dcf),
	.w7(32'hb8282de4),
	.w8(32'h392b3d95),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e98120),
	.w1(32'h384426ae),
	.w2(32'h38de1bcd),
	.w3(32'hb91c0569),
	.w4(32'hb8760023),
	.w5(32'hb782b443),
	.w6(32'hb9199718),
	.w7(32'hb8b554b9),
	.w8(32'hb6896cd1),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb794c94f),
	.w1(32'hb90545c6),
	.w2(32'hb8df544d),
	.w3(32'h38fb0158),
	.w4(32'hb76e2f3a),
	.w5(32'hb819fdb4),
	.w6(32'h395ad0d4),
	.w7(32'h38db4904),
	.w8(32'h39143bc0),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6428a0b),
	.w1(32'hb68bfd78),
	.w2(32'hb7130b5f),
	.w3(32'hb64e77e1),
	.w4(32'hb71fd95c),
	.w5(32'hb6dc3bd0),
	.w6(32'hb5d93dbb),
	.w7(32'hb6da5546),
	.w8(32'hb702d261),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96cbe97),
	.w1(32'hb775fa8c),
	.w2(32'hb8b403ab),
	.w3(32'hb78597c5),
	.w4(32'h393e6b9f),
	.w5(32'h384d236a),
	.w6(32'h38cd9d6c),
	.w7(32'h3930277a),
	.w8(32'h3927296b),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6b0af6e),
	.w1(32'h35522056),
	.w2(32'hb479563c),
	.w3(32'hb67e7421),
	.w4(32'h351093d9),
	.w5(32'h32f94d48),
	.w6(32'hb684b484),
	.w7(32'hb627b43d),
	.w8(32'h349f7bf5),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb721bf03),
	.w1(32'hb6822a9d),
	.w2(32'hb6bd79cc),
	.w3(32'hb688a9e5),
	.w4(32'hb653537f),
	.w5(32'h3698394b),
	.w6(32'hb73bf8f2),
	.w7(32'hb6bc0fdc),
	.w8(32'hb67a9e85),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388cb61c),
	.w1(32'hb9c220a0),
	.w2(32'hb86901a0),
	.w3(32'h38ff51b2),
	.w4(32'hb9c2e8e2),
	.w5(32'hb90044ec),
	.w6(32'h3907d12e),
	.w7(32'hb9a8dc53),
	.w8(32'hb9500646),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ee4c4b),
	.w1(32'hba0b2887),
	.w2(32'h38fc77a0),
	.w3(32'h393c1c0d),
	.w4(32'h3834831c),
	.w5(32'h3a099686),
	.w6(32'h39b674f7),
	.w7(32'hb9216f7a),
	.w8(32'h39dfa3e9),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h378c9bb4),
	.w1(32'hb8b38c31),
	.w2(32'hb7ebc1c8),
	.w3(32'h3830c860),
	.w4(32'hb84f1fe5),
	.w5(32'hb7e92ab5),
	.w6(32'h3915ae42),
	.w7(32'hb7bd516f),
	.w8(32'h362dfbe2),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3932b458),
	.w1(32'hb9c71268),
	.w2(32'hb8fc9b77),
	.w3(32'h39ad79aa),
	.w4(32'hb9348738),
	.w5(32'h379b01fb),
	.w6(32'h39bf0dfc),
	.w7(32'hb8b67d2d),
	.w8(32'hb89ee9c3),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8063917),
	.w1(32'h388a6274),
	.w2(32'h38521bf7),
	.w3(32'h389a0bcc),
	.w4(32'h391403bf),
	.w5(32'hb7369af3),
	.w6(32'hb7db45bb),
	.w7(32'hb7f75c76),
	.w8(32'hb89fdc1e),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb942aaff),
	.w1(32'hb7e59f8e),
	.w2(32'h399540bc),
	.w3(32'hb9162bcd),
	.w4(32'hb7984ad2),
	.w5(32'h38929b16),
	.w6(32'hb9fec5fa),
	.w7(32'hb7ec32a6),
	.w8(32'h39bfb709),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88a0646),
	.w1(32'hb9042b6a),
	.w2(32'h39117023),
	.w3(32'h38665bdd),
	.w4(32'hb888cebf),
	.w5(32'h39418c0a),
	.w6(32'h37b10cc1),
	.w7(32'hb9142460),
	.w8(32'h391ce6ea),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e50c3a),
	.w1(32'h398a1a04),
	.w2(32'h3965cc9c),
	.w3(32'h388484d6),
	.w4(32'h39cee0b0),
	.w5(32'h39edabb7),
	.w6(32'hb86f8509),
	.w7(32'h39766e50),
	.w8(32'h3a09b540),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5a305a3),
	.w1(32'hb6ab4143),
	.w2(32'hb67f967d),
	.w3(32'hb6460236),
	.w4(32'hb6bf30a9),
	.w5(32'hb6e63110),
	.w6(32'hb78f534f),
	.w7(32'hb6015456),
	.w8(32'hb7116655),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7407d13),
	.w1(32'hb8655e49),
	.w2(32'h3906c194),
	.w3(32'hb6f208b1),
	.w4(32'h37e7b621),
	.w5(32'h38dc3116),
	.w6(32'hb7f645bb),
	.w7(32'hb7be19ce),
	.w8(32'h38c5b97d),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5e7fb42),
	.w1(32'h3686fc23),
	.w2(32'h33fb7406),
	.w3(32'hb6b541d7),
	.w4(32'h34dab948),
	.w5(32'hb6385493),
	.w6(32'hb66b9911),
	.w7(32'hb4a85941),
	.w8(32'hb680a5dc),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37a4706f),
	.w1(32'h381ca2b8),
	.w2(32'h37e71d7a),
	.w3(32'h385d6b39),
	.w4(32'h388a185e),
	.w5(32'h372d65cb),
	.w6(32'h388981a7),
	.w7(32'h387f272a),
	.w8(32'h37fe2adb),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a62d69),
	.w1(32'hb8f96237),
	.w2(32'h371132a9),
	.w3(32'h3889df5c),
	.w4(32'hb8f1239d),
	.w5(32'h345f406f),
	.w6(32'h38e2455e),
	.w7(32'hb84a691b),
	.w8(32'h37b3e8b1),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h384f194d),
	.w1(32'hb60d307a),
	.w2(32'h38ccf727),
	.w3(32'h3944da91),
	.w4(32'h3883059d),
	.w5(32'h3911830f),
	.w6(32'h38c8980f),
	.w7(32'h3826c66c),
	.w8(32'h391263c5),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5b3531a),
	.w1(32'h36585865),
	.w2(32'h35dbb91a),
	.w3(32'hb6967a1d),
	.w4(32'h3622bc4f),
	.w5(32'h354c24c2),
	.w6(32'h346e4fe8),
	.w7(32'h362bcfd2),
	.w8(32'hb5b81860),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb475e05d),
	.w1(32'h35f09011),
	.w2(32'h367c4041),
	.w3(32'hb498f709),
	.w4(32'h362b5a5f),
	.w5(32'h35fe6d64),
	.w6(32'h341cfca1),
	.w7(32'h34f58a4f),
	.w8(32'hb5f4aaac),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h380a4d38),
	.w1(32'hb9162138),
	.w2(32'h3768a436),
	.w3(32'h3923c181),
	.w4(32'hb8bdefba),
	.w5(32'h3904d402),
	.w6(32'h39112777),
	.w7(32'h38108924),
	.w8(32'h3829e08a),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9741348),
	.w1(32'hb9a3da38),
	.w2(32'h3875cc26),
	.w3(32'h392ee852),
	.w4(32'hb95b0326),
	.w5(32'hb893484a),
	.w6(32'hb92f52d3),
	.w7(32'hb995ba85),
	.w8(32'hb8c03c6c),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9596801),
	.w1(32'hb906b097),
	.w2(32'h39b16f92),
	.w3(32'hb70985a4),
	.w4(32'hb8fc8d4e),
	.w5(32'h39cbdfc0),
	.w6(32'hb850343c),
	.w7(32'hb9a88705),
	.w8(32'h3941ab50),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h377a6884),
	.w1(32'h36b24c1b),
	.w2(32'hb7d3680d),
	.w3(32'h392b1b33),
	.w4(32'h384ff25a),
	.w5(32'h38da6d11),
	.w6(32'h378b3f1d),
	.w7(32'h3853e941),
	.w8(32'h391f060c),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a7a36b),
	.w1(32'h39ed76df),
	.w2(32'h39e747d9),
	.w3(32'hb66f91d9),
	.w4(32'h39fc9de1),
	.w5(32'h3a12d635),
	.w6(32'hb9946c91),
	.w7(32'h39c7b56b),
	.w8(32'h3a4cf6a1),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b3d194),
	.w1(32'hb9dea1d9),
	.w2(32'h39a48b80),
	.w3(32'h39cf202c),
	.w4(32'hb9ba4ac6),
	.w5(32'hb93ac81f),
	.w6(32'h39c85d0a),
	.w7(32'hb9ae5161),
	.w8(32'hb906d8e4),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96e1ac9),
	.w1(32'h37afd210),
	.w2(32'h39170380),
	.w3(32'hb8c93b7f),
	.w4(32'h39061d6f),
	.w5(32'h390d2a8e),
	.w6(32'hb88f89cf),
	.w7(32'h3805b606),
	.w8(32'h38193028),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h354657ae),
	.w1(32'hb5daf8e5),
	.w2(32'hb63859d3),
	.w3(32'hb64c7f15),
	.w4(32'hb6aa47e5),
	.w5(32'h34cff745),
	.w6(32'hb64b1c2d),
	.w7(32'h363b0794),
	.w8(32'hb622ffca),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb59e5ea5),
	.w1(32'h36a3a999),
	.w2(32'h370f331d),
	.w3(32'hb52d4b15),
	.w4(32'h3650cf10),
	.w5(32'h3700e09c),
	.w6(32'h369f2383),
	.w7(32'h3696859e),
	.w8(32'h37096a45),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb647baa2),
	.w1(32'h36531b6f),
	.w2(32'hb51de184),
	.w3(32'hb69eb161),
	.w4(32'h359e42da),
	.w5(32'hb5e2e483),
	.w6(32'hb61d2192),
	.w7(32'h3589714d),
	.w8(32'hb4d40575),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9edab1d),
	.w1(32'h3809ecbf),
	.w2(32'h38793d93),
	.w3(32'hb9274848),
	.w4(32'h38f2a6f3),
	.w5(32'h360f4406),
	.w6(32'hb90c732b),
	.w7(32'h36a930a6),
	.w8(32'h38170791),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92096db),
	.w1(32'hb955d269),
	.w2(32'h381c41e8),
	.w3(32'hb8a36270),
	.w4(32'hb9195935),
	.w5(32'h38d89d32),
	.w6(32'hb830f723),
	.w7(32'hb9287748),
	.w8(32'h392baf7a),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39674d57),
	.w1(32'hb9b4bd8f),
	.w2(32'h386db76b),
	.w3(32'h39a7a123),
	.w4(32'hb9904f06),
	.w5(32'hb8b752e4),
	.w6(32'h39d50bf1),
	.w7(32'hb9013bb6),
	.w8(32'hb77e6764),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36ee7f75),
	.w1(32'hb8e109d5),
	.w2(32'hb887986f),
	.w3(32'h38e51b32),
	.w4(32'hb87f9218),
	.w5(32'h371b7080),
	.w6(32'h38e445f0),
	.w7(32'hb56d5956),
	.w8(32'h378fbe45),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98c75d0),
	.w1(32'hb901b2af),
	.w2(32'hb880bdd1),
	.w3(32'hb80fcdfa),
	.w4(32'h35db2cce),
	.w5(32'hb7221b98),
	.w6(32'hb82b310d),
	.w7(32'hb80ebc9a),
	.w8(32'h392b8312),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90496e2),
	.w1(32'hb7e9e061),
	.w2(32'h392b4441),
	.w3(32'hb8849d1a),
	.w4(32'h386ce5f5),
	.w5(32'h392c3298),
	.w6(32'hb83218b6),
	.w7(32'hb8097451),
	.w8(32'h383ff5f1),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb635b16d),
	.w1(32'h36493da8),
	.w2(32'hb4da70af),
	.w3(32'hb69c0078),
	.w4(32'h355e2cae),
	.w5(32'hb62dd944),
	.w6(32'hb66731a2),
	.w7(32'h359d748a),
	.w8(32'hb61cac10),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c6451f),
	.w1(32'h36834d82),
	.w2(32'h390bca14),
	.w3(32'hb7733fa4),
	.w4(32'h37b001f2),
	.w5(32'h38e506b9),
	.w6(32'h389e6c95),
	.w7(32'h37e897ed),
	.w8(32'hb895322e),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb51e2ba7),
	.w1(32'h367c9645),
	.w2(32'hb5b7ffc2),
	.w3(32'hb711fb45),
	.w4(32'hb5b8cfd4),
	.w5(32'hb6bf6860),
	.w6(32'hb6ff8383),
	.w7(32'h3601a865),
	.w8(32'hb6e555e5),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb986b9b6),
	.w1(32'hb72a68b0),
	.w2(32'h38658c55),
	.w3(32'hb8b44468),
	.w4(32'h37ba8eb8),
	.w5(32'h392f0571),
	.w6(32'hb885cc0e),
	.w7(32'h37c6c729),
	.w8(32'h39bf5c54),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3968f355),
	.w1(32'hb9fd3874),
	.w2(32'h38688f81),
	.w3(32'h3994c2fd),
	.w4(32'hb9f2f0c7),
	.w5(32'h3785db62),
	.w6(32'h39c544e1),
	.w7(32'hb9a09dde),
	.w8(32'hb8fd1f64),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38eb7932),
	.w1(32'hb9a7825f),
	.w2(32'h3720684d),
	.w3(32'h39aa0eeb),
	.w4(32'hb9268281),
	.w5(32'h38665162),
	.w6(32'h39a5840f),
	.w7(32'hb8e0855c),
	.w8(32'h38272c8a),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37a1f084),
	.w1(32'hb84364e7),
	.w2(32'hb7d1ecb0),
	.w3(32'h3803a9dd),
	.w4(32'hb850c346),
	.w5(32'hb80ce117),
	.w6(32'h386aad50),
	.w7(32'hb823b4d2),
	.w8(32'hb810109e),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397e53ed),
	.w1(32'hb9ef23ea),
	.w2(32'h378f8903),
	.w3(32'h3a057076),
	.w4(32'hb91eb962),
	.w5(32'h38dfc805),
	.w6(32'h3a196b64),
	.w7(32'hb8a641fa),
	.w8(32'h37f2025e),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c41fee),
	.w1(32'hb8c48b41),
	.w2(32'hb830a558),
	.w3(32'h38a3085b),
	.w4(32'h35efb530),
	.w5(32'h387e2049),
	.w6(32'h3796f82e),
	.w7(32'hb7a7f711),
	.w8(32'h38942b65),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f0af23),
	.w1(32'hb95550e4),
	.w2(32'h369238aa),
	.w3(32'h38e7bfea),
	.w4(32'hb864d97b),
	.w5(32'h394e022b),
	.w6(32'h39089e74),
	.w7(32'h390d12e4),
	.w8(32'h3a07ee51),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35c39658),
	.w1(32'hb5495463),
	.w2(32'hb6a78939),
	.w3(32'h367dd2fa),
	.w4(32'h3610e01f),
	.w5(32'hb6570867),
	.w6(32'hb5ae7b11),
	.w7(32'hb49f6a94),
	.w8(32'hb6752779),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb705f905),
	.w1(32'hb6723b69),
	.w2(32'h36b0866b),
	.w3(32'hb6de9d70),
	.w4(32'hb687d519),
	.w5(32'hb5a704ab),
	.w6(32'hb67812a4),
	.w7(32'h36088a68),
	.w8(32'hb52f2443),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bb3ad2),
	.w1(32'hba26ce9b),
	.w2(32'hb863b6e2),
	.w3(32'hb90668ea),
	.w4(32'hb9a57e2f),
	.w5(32'h3858c80c),
	.w6(32'h399b87be),
	.w7(32'hb8c4d40a),
	.w8(32'h3925cdc7),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d0c0fc),
	.w1(32'hb991294d),
	.w2(32'h38c9836e),
	.w3(32'h39c26226),
	.w4(32'h3914c534),
	.w5(32'h3a0c6999),
	.w6(32'h389b2f52),
	.w7(32'hb6aad657),
	.w8(32'h38559437),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h384375f0),
	.w1(32'hb9e971ac),
	.w2(32'hb541c297),
	.w3(32'h39a343f7),
	.w4(32'hb9b892ac),
	.w5(32'h3760b6b6),
	.w6(32'h39748e92),
	.w7(32'hb90c5003),
	.w8(32'h37d5a51b),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba195599),
	.w1(32'h392a5d44),
	.w2(32'h38f9f487),
	.w3(32'hb7b13266),
	.w4(32'h39dc8c97),
	.w5(32'h39152ddc),
	.w6(32'hb8a0efb7),
	.w7(32'h38d52921),
	.w8(32'h39504fbd),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3742e3bf),
	.w1(32'h3676d974),
	.w2(32'hb7bd7409),
	.w3(32'h37baaa82),
	.w4(32'hb6d6550f),
	.w5(32'hb7bd9322),
	.w6(32'h379d45d3),
	.w7(32'h373094d4),
	.w8(32'hb74417bf),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5c26f2e),
	.w1(32'h37f7e12a),
	.w2(32'h3662385f),
	.w3(32'hb844c45f),
	.w4(32'h369cb186),
	.w5(32'h3634d2fc),
	.w6(32'h3800a93c),
	.w7(32'h37ae9a53),
	.w8(32'h35ce1102),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba97b61e),
	.w1(32'hb98cb953),
	.w2(32'h3a0286cc),
	.w3(32'hb9c805bb),
	.w4(32'h384c0b48),
	.w5(32'h3a08752b),
	.w6(32'hb89f4a05),
	.w7(32'hb9a0ae64),
	.w8(32'h39ae41b8),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c8a4f3),
	.w1(32'h39a3ca89),
	.w2(32'h398c3a59),
	.w3(32'hb96356d5),
	.w4(32'h39a03147),
	.w5(32'h3a0efb9a),
	.w6(32'hb951002c),
	.w7(32'h397163ed),
	.w8(32'h3a47fe85),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0cbb46),
	.w1(32'hb93010c9),
	.w2(32'h39bdd354),
	.w3(32'hb95e26b5),
	.w4(32'hb85e103a),
	.w5(32'h39d79887),
	.w6(32'hb8983d53),
	.w7(32'hb9b6023d),
	.w8(32'h39e75373),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e90260),
	.w1(32'hb9bec22c),
	.w2(32'hb8d873ae),
	.w3(32'h39782021),
	.w4(32'hb9931597),
	.w5(32'hb8c05565),
	.w6(32'h39a1b555),
	.w7(32'hb96b6c95),
	.w8(32'hb912c7e5),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d7021c),
	.w1(32'hb9985b20),
	.w2(32'h38d7f478),
	.w3(32'h3a24a54e),
	.w4(32'hb94fc866),
	.w5(32'hb73f6ba8),
	.w6(32'h3a2ceba0),
	.w7(32'hb834c545),
	.w8(32'h37dde351),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb3593f4e),
	.w1(32'hb5d4fc08),
	.w2(32'hb5879893),
	.w3(32'hb3cf671e),
	.w4(32'h33c8b8d7),
	.w5(32'h347affd8),
	.w6(32'hb615c947),
	.w7(32'hb4c07c5d),
	.w8(32'hb5584ede),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb61a1c66),
	.w1(32'h360b4999),
	.w2(32'hb6249a88),
	.w3(32'hb649e5ef),
	.w4(32'h3611097a),
	.w5(32'hb5c47544),
	.w6(32'hb691f168),
	.w7(32'hb609a1df),
	.w8(32'hb6a70199),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98aa1d6),
	.w1(32'hb8db2166),
	.w2(32'hb8b39456),
	.w3(32'hb8d3402f),
	.w4(32'h36690242),
	.w5(32'hb8381cf9),
	.w6(32'h37a5e214),
	.w7(32'h387410ec),
	.w8(32'h3821f542),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb688d8e2),
	.w1(32'h35feb621),
	.w2(32'hb5f9a326),
	.w3(32'hb6cfb74b),
	.w4(32'hb5f1c1d8),
	.w5(32'hb640c27b),
	.w6(32'hb6c74966),
	.w7(32'hb4c15af5),
	.w8(32'hb5fd9541),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb939c4ad),
	.w1(32'h38f229e6),
	.w2(32'h389be895),
	.w3(32'hb8b5710b),
	.w4(32'h391af199),
	.w5(32'h38502092),
	.w6(32'hb81f9d9a),
	.w7(32'h389d94e6),
	.w8(32'h3863d7a6),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90a8e4d),
	.w1(32'hb92e8802),
	.w2(32'h3913f889),
	.w3(32'h37117fe5),
	.w4(32'hb8a640bd),
	.w5(32'h399e0c37),
	.w6(32'h3907a432),
	.w7(32'hb775fb0e),
	.w8(32'h3997b0b0),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h380179f3),
	.w1(32'hb9901dac),
	.w2(32'hb89074d1),
	.w3(32'h3977e61a),
	.w4(32'hb76ac21e),
	.w5(32'h39235737),
	.w6(32'h39827c5b),
	.w7(32'hb8921179),
	.w8(32'hb883a4e0),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb64a9495),
	.w1(32'hb5beedb8),
	.w2(32'hb519b6a8),
	.w3(32'hb73b0bee),
	.w4(32'hb6ac1d6f),
	.w5(32'hb6f57ef6),
	.w6(32'hb5972825),
	.w7(32'hb56a8645),
	.w8(32'hb6d44171),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4b0e9f),
	.w1(32'hb949cb05),
	.w2(32'h3a0000af),
	.w3(32'hb9917643),
	.w4(32'h392032df),
	.w5(32'h3a69e5c0),
	.w6(32'hb93695a7),
	.w7(32'hb9de65a1),
	.w8(32'h3a3e24c1),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93f0610),
	.w1(32'h38969c46),
	.w2(32'h38811300),
	.w3(32'hb8bfa219),
	.w4(32'h38fb5592),
	.w5(32'h394f982b),
	.w6(32'hb8f0bd4e),
	.w7(32'h3885f468),
	.w8(32'h39846e4b),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6719133),
	.w1(32'h359490d4),
	.w2(32'hb5eefb1a),
	.w3(32'hb73fe4f8),
	.w4(32'hb65fd684),
	.w5(32'hb6898849),
	.w6(32'hb619944b),
	.w7(32'h360ac46d),
	.w8(32'hb6c2e706),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b100f7),
	.w1(32'h38b5dba0),
	.w2(32'h38c41698),
	.w3(32'hb9120ddb),
	.w4(32'h39149572),
	.w5(32'h396bacb3),
	.w6(32'hb882b14d),
	.w7(32'h388184bc),
	.w8(32'h39b1f09d),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6880b5d),
	.w1(32'hb67dcfe5),
	.w2(32'hb5d1cbd8),
	.w3(32'hb69cd6bc),
	.w4(32'hb6965095),
	.w5(32'hb64f43e7),
	.w6(32'hb607a6ce),
	.w7(32'hb5c2a31a),
	.w8(32'hb5e5a650),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb644d09a),
	.w1(32'h37069cd9),
	.w2(32'h37ea20c3),
	.w3(32'hb72532e4),
	.w4(32'h369b2ddc),
	.w5(32'h3754c086),
	.w6(32'hb6649646),
	.w7(32'h36fdf5d8),
	.w8(32'h37aa200d),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb66fead8),
	.w1(32'hb5d90aa3),
	.w2(32'h3491ea9a),
	.w3(32'hb66566b1),
	.w4(32'hb2d8865e),
	.w5(32'h33d6b4ce),
	.w6(32'hb5f224ee),
	.w7(32'hb5d3fac7),
	.w8(32'hb628fc02),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6d35e2a),
	.w1(32'hb7007561),
	.w2(32'hb6afa47f),
	.w3(32'hb6f0ffb6),
	.w4(32'hb709aa47),
	.w5(32'hb6718251),
	.w6(32'hb6b8c574),
	.w7(32'hb5f6f45c),
	.w8(32'hb5a5fe13),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8769a17),
	.w1(32'hb967eda7),
	.w2(32'hb864b8b1),
	.w3(32'h38bb7834),
	.w4(32'hb8e44d08),
	.w5(32'h386d2f1d),
	.w6(32'h38da3cc4),
	.w7(32'hb8b1cf6c),
	.w8(32'hb8309f3b),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h373e2a41),
	.w1(32'h397eca8e),
	.w2(32'h395b0733),
	.w3(32'h392fde4d),
	.w4(32'h39b7fd54),
	.w5(32'h39917363),
	.w6(32'hb914a9ee),
	.w7(32'h391487d8),
	.w8(32'h39480b9a),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb96d7c14),
	.w1(32'h389e7205),
	.w2(32'h37be5a3a),
	.w3(32'hb85d9c81),
	.w4(32'h39042c3b),
	.w5(32'h392a0db7),
	.w6(32'hb90a8a09),
	.w7(32'h38202d7c),
	.w8(32'h396bcf16),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97711f8),
	.w1(32'h390bb6ec),
	.w2(32'h38b9b9c9),
	.w3(32'hb7557905),
	.w4(32'h3998791d),
	.w5(32'h392ec0fc),
	.w6(32'hb90b25a1),
	.w7(32'h391c9538),
	.w8(32'h398f10c6),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6b2cebd),
	.w1(32'hb77f4d36),
	.w2(32'hb65f5bba),
	.w3(32'hb7003900),
	.w4(32'hb7732059),
	.w5(32'hb5f24642),
	.w6(32'hb6c53dd6),
	.w7(32'hb74d1b5c),
	.w8(32'hb6e47fe4),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7cc0093),
	.w1(32'h37eefe02),
	.w2(32'hb521c9a4),
	.w3(32'hb7416236),
	.w4(32'h3793d747),
	.w5(32'hb6fe145f),
	.w6(32'hb6987c8d),
	.w7(32'h373f9fd9),
	.w8(32'h367dd093),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb4d4a0df),
	.w1(32'h369c2601),
	.w2(32'h35a9bce3),
	.w3(32'hb62531d8),
	.w4(32'h361d0454),
	.w5(32'h348704e2),
	.w6(32'h3616f23a),
	.w7(32'h36455ce1),
	.w8(32'hb6186cdd),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5450280),
	.w1(32'h366331f3),
	.w2(32'h35a0b53b),
	.w3(32'hb639c30f),
	.w4(32'h35e9757f),
	.w5(32'h3594e324),
	.w6(32'hb58cfcc7),
	.w7(32'h359cd924),
	.w8(32'hb5e9c067),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90bcb7c),
	.w1(32'hb7e03273),
	.w2(32'h390d95a5),
	.w3(32'hb93cda19),
	.w4(32'h389ac1dc),
	.w5(32'h395a350b),
	.w6(32'hb85e27a4),
	.w7(32'h388a666a),
	.w8(32'h39a02dd4),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37284b90),
	.w1(32'h37392618),
	.w2(32'h371b43eb),
	.w3(32'h36f94228),
	.w4(32'h37258b07),
	.w5(32'h36df556d),
	.w6(32'h369bd861),
	.w7(32'h375aca3f),
	.w8(32'h372c5343),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37937607),
	.w1(32'hb7d0a5b1),
	.w2(32'h378265d2),
	.w3(32'h37a70db7),
	.w4(32'hb7a505d9),
	.w5(32'h372e7059),
	.w6(32'h387c6762),
	.w7(32'hb772c0ea),
	.w8(32'h36823184),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a7c5b3),
	.w1(32'hb837b91e),
	.w2(32'h3872de9b),
	.w3(32'h38b85220),
	.w4(32'hb69e1ce7),
	.w5(32'h32e93314),
	.w6(32'h3862e4d5),
	.w7(32'hb81a19be),
	.w8(32'hb754c458),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36384002),
	.w1(32'h36c88717),
	.w2(32'h35cc7a8e),
	.w3(32'h35d9df60),
	.w4(32'h36a63b83),
	.w5(32'h3588b40d),
	.w6(32'h3636de38),
	.w7(32'h36837725),
	.w8(32'hb433c5cc),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8dbef30),
	.w1(32'hb7fb2042),
	.w2(32'h365a6e21),
	.w3(32'hb864d688),
	.w4(32'h384602bf),
	.w5(32'h3890cf51),
	.w6(32'hb8b16b35),
	.w7(32'h37f9e596),
	.w8(32'h3909eea9),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7a16a70),
	.w1(32'h37444cc9),
	.w2(32'hb690f84d),
	.w3(32'hb75aa15b),
	.w4(32'h36c5717c),
	.w5(32'hb6e1e036),
	.w6(32'hb703d76b),
	.w7(32'hb449d13d),
	.w8(32'hb6df19d2),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb815b4b2),
	.w1(32'h39809e1c),
	.w2(32'h39e60f41),
	.w3(32'hb87964c6),
	.w4(32'h39aae069),
	.w5(32'h39bb613d),
	.w6(32'hb9b871c8),
	.w7(32'h38a5c0f8),
	.w8(32'h39f3c1cb),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb68bf166),
	.w1(32'hbafbc548),
	.w2(32'hbb67a60d),
	.w3(32'hb64f33c9),
	.w4(32'h399e49ce),
	.w5(32'hbafdcaf3),
	.w6(32'hba88f6dc),
	.w7(32'hbb62ed39),
	.w8(32'hbac37f6c),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae7de54),
	.w1(32'hba2f3ded),
	.w2(32'h3a9a8ddc),
	.w3(32'hba6e249c),
	.w4(32'h39746122),
	.w5(32'h39da5704),
	.w6(32'hb9be9386),
	.w7(32'h3a5da1d7),
	.w8(32'h3a0ac417),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule