module layer_10_featuremap_85(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b42ac69),
	.w1(32'hbc157985),
	.w2(32'hbb16854f),
	.w3(32'hbacb03e9),
	.w4(32'h3b4fb295),
	.w5(32'h3b295177),
	.w6(32'h3ca41ecc),
	.w7(32'h3a676a03),
	.w8(32'h3ad80d8a),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d26a2e3),
	.w1(32'h3b649be6),
	.w2(32'hbb18f90a),
	.w3(32'h3b091baf),
	.w4(32'hbb9a3072),
	.w5(32'h3abdcf7a),
	.w6(32'h3b33aadc),
	.w7(32'h3ae0a8b4),
	.w8(32'h3b7ff2c9),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b401afb),
	.w1(32'h3b182fd1),
	.w2(32'h3a98714d),
	.w3(32'hba0c555f),
	.w4(32'h3c8fa7c9),
	.w5(32'h3c191f6c),
	.w6(32'hba12bf2e),
	.w7(32'hba1c582d),
	.w8(32'h3ae3470a),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab35884),
	.w1(32'h3b04e1a0),
	.w2(32'h3a67a4c9),
	.w3(32'h3ba20dec),
	.w4(32'h3c036955),
	.w5(32'h3b79b951),
	.w6(32'h3922d65a),
	.w7(32'h3afed752),
	.w8(32'hbbbb4e82),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb685b6a),
	.w1(32'hbb53d1c5),
	.w2(32'h38d9c8ca),
	.w3(32'hbb82d87b),
	.w4(32'h3a2bec17),
	.w5(32'hbb160f2e),
	.w6(32'hbb5a8175),
	.w7(32'hb9c1a38a),
	.w8(32'h3c85b54b),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb63be77),
	.w1(32'hbb660e99),
	.w2(32'h3b124da1),
	.w3(32'hbb881f79),
	.w4(32'h3a8ac4c5),
	.w5(32'h3bd6e415),
	.w6(32'h3b91f80d),
	.w7(32'hba95a3e5),
	.w8(32'h3baed6f2),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e3cde8),
	.w1(32'h3b4a8de8),
	.w2(32'hbb08f4da),
	.w3(32'hbb4aea47),
	.w4(32'hbc593034),
	.w5(32'hbb04eb54),
	.w6(32'hbaae7894),
	.w7(32'hbb803359),
	.w8(32'hbb910b51),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd9d2c8),
	.w1(32'hba6bb42d),
	.w2(32'h3b5f0d4e),
	.w3(32'hbba411cf),
	.w4(32'h3a6e7a5e),
	.w5(32'h39ae87ab),
	.w6(32'hbbf457ce),
	.w7(32'hbbb41ca2),
	.w8(32'hbacffd20),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c433226),
	.w1(32'hbcb9f1c1),
	.w2(32'h3b95385f),
	.w3(32'h3acfcc02),
	.w4(32'h3b2b1aba),
	.w5(32'hba1825c8),
	.w6(32'hbbb37706),
	.w7(32'hbb28c890),
	.w8(32'hb9a1571d),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8241f9),
	.w1(32'h39d363a4),
	.w2(32'h3c059e06),
	.w3(32'hb9d267f8),
	.w4(32'h3af9aeb9),
	.w5(32'h38b5c178),
	.w6(32'h3b32d682),
	.w7(32'h3ba161ad),
	.w8(32'h3b33762e),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc2f122),
	.w1(32'h3a3857c4),
	.w2(32'hbb072a2c),
	.w3(32'hba811e9e),
	.w4(32'hbc32c5e0),
	.w5(32'h3cb51f47),
	.w6(32'h3ac3b07b),
	.w7(32'hbb21837b),
	.w8(32'hbb04d1cb),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cad21e0),
	.w1(32'hbb47699f),
	.w2(32'h38ce48c2),
	.w3(32'h39fa8793),
	.w4(32'hbbccddde),
	.w5(32'hb7c53dd0),
	.w6(32'hbaa92c59),
	.w7(32'hba03ec83),
	.w8(32'hba190523),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2e2bb2),
	.w1(32'hbab3e2a5),
	.w2(32'h3ba33c24),
	.w3(32'hbb9ce84b),
	.w4(32'hbabecb90),
	.w5(32'h3a3be967),
	.w6(32'hbb38cd4f),
	.w7(32'h3b96cd23),
	.w8(32'h39a87a87),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca06ff9),
	.w1(32'h3aac3ffd),
	.w2(32'hbad9fc24),
	.w3(32'hba122030),
	.w4(32'h395b20cb),
	.w5(32'h3aab271c),
	.w6(32'h3b2da4f8),
	.w7(32'hbca622fc),
	.w8(32'h39805eef),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafdb19e),
	.w1(32'hba6e0970),
	.w2(32'hbb279087),
	.w3(32'hbaf5ca6e),
	.w4(32'h3b675cbf),
	.w5(32'h3b935243),
	.w6(32'hba2cc876),
	.w7(32'h3b014050),
	.w8(32'hb9ff076b),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aee2873),
	.w1(32'hbacd0704),
	.w2(32'h3a89aa45),
	.w3(32'hbc0bed8f),
	.w4(32'h3a64824e),
	.w5(32'h3b08d746),
	.w6(32'h3b8cebbd),
	.w7(32'hbb185c1f),
	.w8(32'hbc7e3a72),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba40b423),
	.w1(32'hbc6b4450),
	.w2(32'h3b5ebe36),
	.w3(32'hbadcb861),
	.w4(32'hb8535ad1),
	.w5(32'h3c0b7bd7),
	.w6(32'h3b36ab79),
	.w7(32'hbb77f005),
	.w8(32'hba87d7ce),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5f113b),
	.w1(32'h3ce51307),
	.w2(32'h3cc9a6f1),
	.w3(32'h3b0bbdec),
	.w4(32'hba64c901),
	.w5(32'h3ab324cd),
	.w6(32'h3b39ddd4),
	.w7(32'h3bc7e631),
	.w8(32'hba704249),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb278c82),
	.w1(32'h3c1d9dba),
	.w2(32'h3b3b2aa6),
	.w3(32'h3adff387),
	.w4(32'hba637124),
	.w5(32'h3b9b0e41),
	.w6(32'hbb1d79f5),
	.w7(32'hbb8d7a3e),
	.w8(32'h3a1b6c65),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c99bf73),
	.w1(32'hbad68d8e),
	.w2(32'hbae8fb90),
	.w3(32'h3a98dd3b),
	.w4(32'hbbc5bfbb),
	.w5(32'h3a45e953),
	.w6(32'hbb15c610),
	.w7(32'hba096956),
	.w8(32'hba25fa7d),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaa06bc),
	.w1(32'hba54894e),
	.w2(32'hbc247bfc),
	.w3(32'h3979ec48),
	.w4(32'h3ab61b99),
	.w5(32'hbb6db9cb),
	.w6(32'hbbca81ab),
	.w7(32'hba635677),
	.w8(32'h3a9c952c),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc08dae3),
	.w1(32'hbab14d43),
	.w2(32'h3bc8baf2),
	.w3(32'h39c52285),
	.w4(32'hbb514479),
	.w5(32'h38d9f912),
	.w6(32'hba83f17e),
	.w7(32'h39925d58),
	.w8(32'hbb5dfc60),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3949bfc6),
	.w1(32'hb913ea36),
	.w2(32'hbc08fee3),
	.w3(32'h39e9fa3b),
	.w4(32'hbb66da92),
	.w5(32'h3cb22f3c),
	.w6(32'hbb2c0eff),
	.w7(32'hbba0eaa3),
	.w8(32'hbb0da3ab),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb18a82f),
	.w1(32'hbb2abff5),
	.w2(32'hba828eb0),
	.w3(32'hba0f0735),
	.w4(32'hba74ecc0),
	.w5(32'h3afab2b6),
	.w6(32'hbb7af23b),
	.w7(32'hbb238fb7),
	.w8(32'h38994360),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa05d2a),
	.w1(32'h39834b52),
	.w2(32'hb9d7ba20),
	.w3(32'hbae81d83),
	.w4(32'hb9c32ecf),
	.w5(32'hbaf17159),
	.w6(32'h3923fa22),
	.w7(32'h3ae5ed36),
	.w8(32'hba6dc2b6),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be6ef03),
	.w1(32'hb9a6c317),
	.w2(32'hb992ca3e),
	.w3(32'h3bccac82),
	.w4(32'hbb19ff56),
	.w5(32'hbb1c5379),
	.w6(32'hbbf06945),
	.w7(32'h38d110b5),
	.w8(32'h3b8cd0f2),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4a35b5),
	.w1(32'hbb191ac6),
	.w2(32'h38820d7c),
	.w3(32'hb9ba66e5),
	.w4(32'hb99903fa),
	.w5(32'h3b2017e0),
	.w6(32'h3bafdde7),
	.w7(32'hbb4a5ec4),
	.w8(32'h3a18c0ba),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adaf8b7),
	.w1(32'hbba8b953),
	.w2(32'h3a56cb80),
	.w3(32'h3b6cd6ee),
	.w4(32'hbb5702e2),
	.w5(32'h3ccb74eb),
	.w6(32'h3adee1d4),
	.w7(32'hbc1c04af),
	.w8(32'hbab41461),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aab2905),
	.w1(32'h39c151ab),
	.w2(32'hbc9336e5),
	.w3(32'hbb9fa55d),
	.w4(32'h3a633402),
	.w5(32'hbacc7d6c),
	.w6(32'h3a552f79),
	.w7(32'hba1399e1),
	.w8(32'h3b557518),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b528a52),
	.w1(32'h3acec092),
	.w2(32'h398958d8),
	.w3(32'hb9c4006c),
	.w4(32'hbc8be754),
	.w5(32'hb95eca54),
	.w6(32'h3a016bd7),
	.w7(32'h3b0e3555),
	.w8(32'hba91e100),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a321711),
	.w1(32'h3a15dac1),
	.w2(32'h3ac8efe3),
	.w3(32'h3af0ef18),
	.w4(32'h3af1498b),
	.w5(32'h3a734625),
	.w6(32'h3aa91577),
	.w7(32'h3a4034cb),
	.w8(32'h3b0f50fd),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d56616),
	.w1(32'hba0261c2),
	.w2(32'h395d21de),
	.w3(32'h3b1a29c2),
	.w4(32'hb85f1138),
	.w5(32'h3a1a76f3),
	.w6(32'h398e6f84),
	.w7(32'hba3434a2),
	.w8(32'h39e8830a),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4203c5),
	.w1(32'hbadcf842),
	.w2(32'h3a33814b),
	.w3(32'h3aad92ca),
	.w4(32'h3b0ff90a),
	.w5(32'h3b00d9ab),
	.w6(32'h3a4a65c5),
	.w7(32'h3aaf91a4),
	.w8(32'hba392b44),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae1f385),
	.w1(32'h3c014138),
	.w2(32'hbbb09f60),
	.w3(32'h3aff1fbd),
	.w4(32'h3a33e421),
	.w5(32'hbb09697b),
	.w6(32'hb71240b7),
	.w7(32'h3b457809),
	.w8(32'h3909bca4),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5d4ae4),
	.w1(32'h3ad90337),
	.w2(32'hbaf2e29e),
	.w3(32'h3b41e29b),
	.w4(32'h3a139a06),
	.w5(32'h3a2516d0),
	.w6(32'hb8d29777),
	.w7(32'h3aa68b54),
	.w8(32'hbc3db92d),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7c58f4),
	.w1(32'h3adc68d1),
	.w2(32'h39b41a73),
	.w3(32'h3b00f90c),
	.w4(32'hbb852c36),
	.w5(32'h3afe9042),
	.w6(32'h3cab7f58),
	.w7(32'h3984819c),
	.w8(32'hbb16c056),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb83767a7),
	.w1(32'h3b2f6487),
	.w2(32'hbb6b2820),
	.w3(32'hbbd8f7da),
	.w4(32'hbbcf0f2f),
	.w5(32'h3cb1f3d3),
	.w6(32'h3abfd6fe),
	.w7(32'hba02c70d),
	.w8(32'h39cca85a),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5617d0),
	.w1(32'h39505dc5),
	.w2(32'h3b0cf78e),
	.w3(32'h38ac177f),
	.w4(32'hbb919f3a),
	.w5(32'hbaa35939),
	.w6(32'hb8c66702),
	.w7(32'hbad83cda),
	.w8(32'hb8aa653e),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2a3c4c),
	.w1(32'hba24199a),
	.w2(32'hbb69fd76),
	.w3(32'h38e83f43),
	.w4(32'h3a737d8c),
	.w5(32'hb9f2de08),
	.w6(32'h399dcce1),
	.w7(32'h3a19ecc1),
	.w8(32'hba6128d6),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0242cf),
	.w1(32'h3a001a91),
	.w2(32'h3a0761e0),
	.w3(32'h3a5bd042),
	.w4(32'hbc522173),
	.w5(32'hba1f0da6),
	.w6(32'hbcb34175),
	.w7(32'h3918cdbd),
	.w8(32'hbb32f3c8),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37f62ceb),
	.w1(32'hb9ae31fa),
	.w2(32'h3aaeaa8c),
	.w3(32'hba2c6c7f),
	.w4(32'h3a1a7c1b),
	.w5(32'h3aad7e46),
	.w6(32'h383a2031),
	.w7(32'h3a2d5f29),
	.w8(32'h39084027),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1a4395),
	.w1(32'h3a14f2fa),
	.w2(32'h3b484531),
	.w3(32'h3aa62b13),
	.w4(32'h3d10d9cf),
	.w5(32'hbb928716),
	.w6(32'h3a99ea21),
	.w7(32'hbaa40860),
	.w8(32'hbb5bac6f),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c42c574),
	.w1(32'h3a91b950),
	.w2(32'hbb340ae4),
	.w3(32'hbab2a7a0),
	.w4(32'hbb093ee9),
	.w5(32'hbaaf53e3),
	.w6(32'hb9d43aa1),
	.w7(32'hbb2f1909),
	.w8(32'h3ac26370),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab9fff4),
	.w1(32'h3b064cb9),
	.w2(32'h3a8a40d6),
	.w3(32'h3ac928e7),
	.w4(32'h39855a12),
	.w5(32'h3b3bfce8),
	.w6(32'h3ba7f9ab),
	.w7(32'h3c7417d2),
	.w8(32'h39b8e4fe),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1767fb),
	.w1(32'h3cb53fe3),
	.w2(32'h3b173735),
	.w3(32'h3a3ad269),
	.w4(32'hba349fbd),
	.w5(32'h3ce7cf28),
	.w6(32'h3ac214e7),
	.w7(32'hbb1ef165),
	.w8(32'h3892f8b4),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3553c8),
	.w1(32'h3a8e618e),
	.w2(32'hbad8822b),
	.w3(32'h3b580ef2),
	.w4(32'hbb00bfc2),
	.w5(32'hbc901b7b),
	.w6(32'hbc7b0b9f),
	.w7(32'h3942b93f),
	.w8(32'hbafc36f9),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd495ca),
	.w1(32'h3b049389),
	.w2(32'h3a9cb12a),
	.w3(32'hbc5f0a0b),
	.w4(32'h3b984994),
	.w5(32'hbc114d0d),
	.w6(32'h39f4ee82),
	.w7(32'h3b3420ae),
	.w8(32'h38ee888f),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c564b),
	.w1(32'h3b572e89),
	.w2(32'h3b5f6c79),
	.w3(32'h38fe5d1b),
	.w4(32'hbc117e25),
	.w5(32'h3b84fca0),
	.w6(32'h3b4e082c),
	.w7(32'hb8d321c9),
	.w8(32'hbbdf16ac),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d742ae),
	.w1(32'hbac6e2e6),
	.w2(32'h3b907769),
	.w3(32'hbad6bada),
	.w4(32'hbb099f29),
	.w5(32'h3ae91630),
	.w6(32'h3a3b6a55),
	.w7(32'h3a878e9f),
	.w8(32'hba0f13de),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b029843),
	.w1(32'hb93b4987),
	.w2(32'h39eb661f),
	.w3(32'hbb663e6d),
	.w4(32'h3aa763b0),
	.w5(32'h3a89d4c6),
	.w6(32'hbae09e55),
	.w7(32'h3a35c124),
	.w8(32'hb9d15694),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93a2e6c),
	.w1(32'h3a92b245),
	.w2(32'hbaac56b1),
	.w3(32'h3aa83bdb),
	.w4(32'h3ab656b7),
	.w5(32'h38d66b12),
	.w6(32'hb9c850f7),
	.w7(32'h3adeb390),
	.w8(32'hba0aec7e),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeea02b),
	.w1(32'hbac9e398),
	.w2(32'h3aa492c3),
	.w3(32'hbb53c9a0),
	.w4(32'hbb42c35c),
	.w5(32'hbb286a68),
	.w6(32'hbc45dff9),
	.w7(32'h3ab73314),
	.w8(32'hb9bdf7df),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aef80e2),
	.w1(32'hbacab107),
	.w2(32'hb9c751e0),
	.w3(32'hba612ed1),
	.w4(32'h3abc91b0),
	.w5(32'hba346397),
	.w6(32'h3ab6479e),
	.w7(32'h3ae0d032),
	.w8(32'h3aa853a2),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7be5f3),
	.w1(32'h3b059ee1),
	.w2(32'hb8c12370),
	.w3(32'h3acce3c8),
	.w4(32'h3b064829),
	.w5(32'hbb2a3b62),
	.w6(32'h3ab060f2),
	.w7(32'h3aed97cd),
	.w8(32'hbb198754),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b9caa7),
	.w1(32'h3ab4513a),
	.w2(32'h3b11d79e),
	.w3(32'h3adad4a6),
	.w4(32'hbb70b313),
	.w5(32'h3af3914a),
	.w6(32'h3a9b3aca),
	.w7(32'h3b797c33),
	.w8(32'h3a65fccd),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb81054f9),
	.w1(32'hbb1d1e33),
	.w2(32'hba556486),
	.w3(32'hb9a98976),
	.w4(32'h3b3afc76),
	.w5(32'hbac47e8b),
	.w6(32'h3a491fac),
	.w7(32'h3a2d831b),
	.w8(32'hbb364726),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aee7f13),
	.w1(32'hbab32271),
	.w2(32'h3c06a672),
	.w3(32'hba3bc51e),
	.w4(32'hb91de844),
	.w5(32'h3aa1d96c),
	.w6(32'hbcb1d2c5),
	.w7(32'hbb1a8c88),
	.w8(32'h3b04bc4b),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb39bfd8),
	.w1(32'h3a5fff47),
	.w2(32'hbb7db7e7),
	.w3(32'h3d0fbc88),
	.w4(32'h3862be74),
	.w5(32'h3b43c6f0),
	.w6(32'hb91421c9),
	.w7(32'h3ae31c8c),
	.w8(32'h3d05b341),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bda066d),
	.w1(32'h3ba6503c),
	.w2(32'h39cce5d3),
	.w3(32'h3ac5e854),
	.w4(32'hba280c12),
	.w5(32'h36619223),
	.w6(32'hb9b8c9e2),
	.w7(32'hbae0985d),
	.w8(32'h3932a12c),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9d8807),
	.w1(32'h3b6ffb54),
	.w2(32'h39cb3a41),
	.w3(32'hbbacba6d),
	.w4(32'hbb07b12d),
	.w5(32'h3b3c1362),
	.w6(32'hbb02298b),
	.w7(32'hbae67b84),
	.w8(32'h3bbe05a4),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad5ab53),
	.w1(32'h3a59765d),
	.w2(32'h39fbaef3),
	.w3(32'hb8c54c00),
	.w4(32'h3bbcd5a8),
	.w5(32'h395366dd),
	.w6(32'h3ac5c5f4),
	.w7(32'h3b0470b2),
	.w8(32'hbb02b0a8),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab638a8),
	.w1(32'hb9d3571a),
	.w2(32'hba27d043),
	.w3(32'hbb1f9edc),
	.w4(32'h3ae95b40),
	.w5(32'hbadd9bc3),
	.w6(32'hbb09824c),
	.w7(32'h3abc89a9),
	.w8(32'h3b4702d4),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4aeaa8),
	.w1(32'h3b2b15a9),
	.w2(32'hbb316ef7),
	.w3(32'h3c1528e2),
	.w4(32'hba0665f4),
	.w5(32'hba3e8bf3),
	.w6(32'h3a8a1946),
	.w7(32'hbb6e9bc8),
	.w8(32'h3a4b4ad1),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd4b0d0),
	.w1(32'h3a213005),
	.w2(32'hbafa9536),
	.w3(32'hba6c2375),
	.w4(32'h3b0bdb40),
	.w5(32'hbbcaf445),
	.w6(32'h3c1b6604),
	.w7(32'hba0e1ec4),
	.w8(32'h3aa8364a),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb80ccac),
	.w1(32'hbb0865fb),
	.w2(32'h3adf97cd),
	.w3(32'h3b263481),
	.w4(32'hbb73a1a1),
	.w5(32'h3b1e1e27),
	.w6(32'h3b942e0e),
	.w7(32'h3beaaba2),
	.w8(32'h3b8edb02),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5c1ed4),
	.w1(32'h3b16af5b),
	.w2(32'hba9e2e84),
	.w3(32'h3b5fe5ec),
	.w4(32'h3a82b746),
	.w5(32'hb7d93425),
	.w6(32'hbc15876c),
	.w7(32'h3c5372bc),
	.w8(32'h3bd0659b),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a84e4be),
	.w1(32'hb9960fd9),
	.w2(32'hba68413d),
	.w3(32'h3c093252),
	.w4(32'hbb62fde1),
	.w5(32'hbb3af824),
	.w6(32'hb6a20583),
	.w7(32'h3be84e22),
	.w8(32'h3a4f77a9),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc07b89),
	.w1(32'hbbb381bd),
	.w2(32'h3ccae284),
	.w3(32'hbb6ab685),
	.w4(32'hbac2a9d3),
	.w5(32'hb7d3a4a9),
	.w6(32'h3a902294),
	.w7(32'hbb5934ef),
	.w8(32'h3c8e24c7),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6102e9),
	.w1(32'h397a446d),
	.w2(32'h39abf7e2),
	.w3(32'hbb03f0bf),
	.w4(32'h38bc4474),
	.w5(32'h393ef98a),
	.w6(32'h3b82b7f4),
	.w7(32'hbb878721),
	.w8(32'h3b411349),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab5e842),
	.w1(32'hbb13332d),
	.w2(32'h3b4caff3),
	.w3(32'h3a4a244e),
	.w4(32'hba8ef19f),
	.w5(32'h38d203fd),
	.w6(32'hbaf97447),
	.w7(32'hbb8dec81),
	.w8(32'hbc79e087),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b186b40),
	.w1(32'hbb84b3e9),
	.w2(32'h3b352628),
	.w3(32'h3bd35045),
	.w4(32'hbcad7bd2),
	.w5(32'hbabee966),
	.w6(32'hbc073104),
	.w7(32'hbbedab6d),
	.w8(32'hbaef56c5),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3262fb),
	.w1(32'h3c0a81cc),
	.w2(32'hbaca4473),
	.w3(32'h38a91119),
	.w4(32'h3a2940ce),
	.w5(32'hbaa21d8f),
	.w6(32'h3850aeaa),
	.w7(32'h3be60959),
	.w8(32'h3b06c19c),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc015fa1),
	.w1(32'hb9836db4),
	.w2(32'h3b07b311),
	.w3(32'h3b082c87),
	.w4(32'hba9bd618),
	.w5(32'hba62e037),
	.w6(32'h3b997ed6),
	.w7(32'h3b118817),
	.w8(32'h3a076459),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afb6dd0),
	.w1(32'h394337db),
	.w2(32'h3b28b283),
	.w3(32'hbb6d2528),
	.w4(32'hba91dad8),
	.w5(32'h39f76d98),
	.w6(32'hbc47b6e0),
	.w7(32'hb9986bcd),
	.w8(32'hbb6d243b),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3fd786),
	.w1(32'h3a126457),
	.w2(32'h389ebc59),
	.w3(32'hbaca18cf),
	.w4(32'h3b45b6ba),
	.w5(32'hbbb07f9a),
	.w6(32'h3c814853),
	.w7(32'h3cc0a496),
	.w8(32'h3902f51c),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0b6042),
	.w1(32'hbb08cb2e),
	.w2(32'hb8afcf89),
	.w3(32'h3a42a59d),
	.w4(32'h3b6f821e),
	.w5(32'hba5661d3),
	.w6(32'h3c86e5bd),
	.w7(32'h3ad0670c),
	.w8(32'h3cc66a6c),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba71a063),
	.w1(32'hbac154c6),
	.w2(32'hbb6ecc9f),
	.w3(32'hba970868),
	.w4(32'h3add0c14),
	.w5(32'h3a043755),
	.w6(32'h3b07d2ea),
	.w7(32'hbae11e16),
	.w8(32'hbb8c531a),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb16ed77),
	.w1(32'hba30bb45),
	.w2(32'hbb02bc3f),
	.w3(32'hbb9631e5),
	.w4(32'hb7d31410),
	.w5(32'h3ac363a0),
	.w6(32'h3b575ead),
	.w7(32'hbaa640b6),
	.w8(32'hbb15ba46),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5ebdf9),
	.w1(32'hb986141e),
	.w2(32'hb889abd3),
	.w3(32'h3ad6eb73),
	.w4(32'h39993c02),
	.w5(32'h3acb900e),
	.w6(32'hbac0d523),
	.w7(32'hba5d422b),
	.w8(32'h3ac9762e),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b439a0b),
	.w1(32'h3a04b2c6),
	.w2(32'hbc4ce66c),
	.w3(32'hba96be7a),
	.w4(32'h3b95d20f),
	.w5(32'h3b8ce0f1),
	.w6(32'hb9b32ec2),
	.w7(32'h3ca50a66),
	.w8(32'h376e31d3),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91acbda),
	.w1(32'h3a8cb89a),
	.w2(32'h3b12b65c),
	.w3(32'h3b38c271),
	.w4(32'h3b00c917),
	.w5(32'hbadc90e6),
	.w6(32'h3ac52a66),
	.w7(32'h3b599333),
	.w8(32'hbaec87fd),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafd304f),
	.w1(32'hbaa362a3),
	.w2(32'h3b61b4ef),
	.w3(32'h3b0005dc),
	.w4(32'h3a82a52d),
	.w5(32'hbab6daae),
	.w6(32'hbb7bd649),
	.w7(32'h3b0a365c),
	.w8(32'h3c1efa17),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6ea671),
	.w1(32'h3ab92832),
	.w2(32'h3a65fe38),
	.w3(32'hbbff806c),
	.w4(32'hbaa0c911),
	.w5(32'hbbbcce91),
	.w6(32'hbb407c1f),
	.w7(32'hba2dfdd5),
	.w8(32'h3b49c666),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb47640e),
	.w1(32'h3b9973e0),
	.w2(32'hb9981293),
	.w3(32'hbb7a7253),
	.w4(32'h3a483fba),
	.w5(32'h3b3b9022),
	.w6(32'hbab43cb7),
	.w7(32'hbb1654b5),
	.w8(32'h3b1c081d),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b017cd8),
	.w1(32'hbbcbac22),
	.w2(32'h3c4ac231),
	.w3(32'hb9412eee),
	.w4(32'hbafc2fad),
	.w5(32'hbb366c10),
	.w6(32'hbb5de3b5),
	.w7(32'hba86ad1a),
	.w8(32'h387bd330),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5a144f),
	.w1(32'h3a8a79e6),
	.w2(32'h3a3eb6d2),
	.w3(32'h3b64af9e),
	.w4(32'h399e847e),
	.w5(32'h3bb591b0),
	.w6(32'h3b6d7dbc),
	.w7(32'hbc883617),
	.w8(32'h3c06f3f7),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b45ed1b),
	.w1(32'hbc6c60ad),
	.w2(32'hbbbb049f),
	.w3(32'h3c2921dc),
	.w4(32'h3a13e9f2),
	.w5(32'hbb46feca),
	.w6(32'h3aefb87e),
	.w7(32'hbb0aa104),
	.w8(32'h3b38c7ba),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba52df7f),
	.w1(32'hbb0beb5d),
	.w2(32'h3bbfbb03),
	.w3(32'h388703e4),
	.w4(32'h3b2a5cc3),
	.w5(32'h3c0edbf8),
	.w6(32'hbb40db61),
	.w7(32'h3c9c7349),
	.w8(32'hba9d08a5),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8d70f2),
	.w1(32'h3af38232),
	.w2(32'h3b1898c1),
	.w3(32'hbb32b8c4),
	.w4(32'hbc08e86a),
	.w5(32'h3b3c49fe),
	.w6(32'h39f2bfeb),
	.w7(32'hbba87d05),
	.w8(32'hb9ee482c),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a99d9bd),
	.w1(32'h3abd8554),
	.w2(32'hb8d59ffe),
	.w3(32'hbb226f7c),
	.w4(32'h3a67c598),
	.w5(32'h39876eba),
	.w6(32'h3aa1794e),
	.w7(32'hba1da765),
	.w8(32'h3b2a390e),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad08fc2),
	.w1(32'hbbca1b34),
	.w2(32'hba397a83),
	.w3(32'h392037a6),
	.w4(32'h3b907c7f),
	.w5(32'hbb0c9a88),
	.w6(32'h3c5ae110),
	.w7(32'hbc02277c),
	.w8(32'hbbf151c4),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acf1d83),
	.w1(32'h3afefaa4),
	.w2(32'h3b1da248),
	.w3(32'h3be9c84d),
	.w4(32'h3bb04a25),
	.w5(32'hbc99af77),
	.w6(32'hba88f152),
	.w7(32'hbb3c82ca),
	.w8(32'h3a7f2cbf),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfb322b),
	.w1(32'hbbfd4ce4),
	.w2(32'h3bcdb8fd),
	.w3(32'h3ab1e00b),
	.w4(32'hbbe923c5),
	.w5(32'hb9928960),
	.w6(32'h3b87c729),
	.w7(32'hbb885b1b),
	.w8(32'h3acbacef),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb28be66),
	.w1(32'hbb223f93),
	.w2(32'h3b576436),
	.w3(32'h3b978152),
	.w4(32'hbb6dac16),
	.w5(32'h3a10a4a8),
	.w6(32'hbb306669),
	.w7(32'hb9c72559),
	.w8(32'hbb004b4d),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b27fb32),
	.w1(32'hbcd04870),
	.w2(32'h39a9db6c),
	.w3(32'h3af0bfb4),
	.w4(32'h3ba10c9a),
	.w5(32'hb9ab2efb),
	.w6(32'h38d2250f),
	.w7(32'h3b175ed6),
	.w8(32'hbaacee0f),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba26546e),
	.w1(32'hbbdc967b),
	.w2(32'hba975585),
	.w3(32'h39d771ee),
	.w4(32'hbbb0f214),
	.w5(32'h39006bef),
	.w6(32'h3b3d28fc),
	.w7(32'h3b6bb60e),
	.w8(32'h39fefed7),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b04e5a6),
	.w1(32'hbc3006f6),
	.w2(32'hbb92ed4a),
	.w3(32'hbc65644d),
	.w4(32'h3b940b73),
	.w5(32'hbce38582),
	.w6(32'hbb730786),
	.w7(32'hbaa48b74),
	.w8(32'hb892d662),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb3d1f7),
	.w1(32'hbb3a6fa7),
	.w2(32'hba98efa9),
	.w3(32'h37fe900c),
	.w4(32'h3aacb266),
	.w5(32'h3abb76e9),
	.w6(32'h3a8d3225),
	.w7(32'h3b10b9f7),
	.w8(32'hbb31ac70),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9da03e),
	.w1(32'h3c8c5aa3),
	.w2(32'hbc31296e),
	.w3(32'h3ae8e52e),
	.w4(32'hbb1b577d),
	.w5(32'h3cd9b91c),
	.w6(32'hbb4600e3),
	.w7(32'h3c08b2d8),
	.w8(32'h3c89ac12),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb361352),
	.w1(32'hbc12c9b7),
	.w2(32'hb8ee8159),
	.w3(32'h3b102aba),
	.w4(32'h3b8f4003),
	.w5(32'h3b4009a2),
	.w6(32'hbba30304),
	.w7(32'hbbc559f1),
	.w8(32'h3b87bf1d),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbdb4b2),
	.w1(32'h3ad44851),
	.w2(32'h39ccf60e),
	.w3(32'hbb07af00),
	.w4(32'hbbd174fe),
	.w5(32'hbbeaa608),
	.w6(32'hbafb68e7),
	.w7(32'hbb512e37),
	.w8(32'hbb6b0461),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa4dfe8),
	.w1(32'h3b2be22b),
	.w2(32'h3c8c91f3),
	.w3(32'h3b1c73de),
	.w4(32'hbb0400bd),
	.w5(32'h394a447e),
	.w6(32'h3c39ce1b),
	.w7(32'hba49f5f5),
	.w8(32'hbb077dc7),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aff211b),
	.w1(32'hbb8dba0a),
	.w2(32'hbc6a76ad),
	.w3(32'hbc11cbd8),
	.w4(32'h3b21653f),
	.w5(32'hbb0aad10),
	.w6(32'hbaefb007),
	.w7(32'hbaf92b5c),
	.w8(32'h3c148d2c),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc21e86a),
	.w1(32'h3bd3fd8e),
	.w2(32'hbbec482d),
	.w3(32'hb98cfbe0),
	.w4(32'h3ae35de7),
	.w5(32'hbba88be4),
	.w6(32'hbabd226b),
	.w7(32'hb97c4d06),
	.w8(32'hbb3a2607),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9ede3d),
	.w1(32'hbc0c24a2),
	.w2(32'h3add4126),
	.w3(32'h3a6a1274),
	.w4(32'hbad44553),
	.w5(32'hbc9aa3f9),
	.w6(32'h3b838d4c),
	.w7(32'hbbda4868),
	.w8(32'hbb5c0f46),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a92930a),
	.w1(32'h3b55a873),
	.w2(32'hb919dabe),
	.w3(32'h38f9fa45),
	.w4(32'h39240cca),
	.w5(32'hba8a783c),
	.w6(32'hba7a45ff),
	.w7(32'hbc179d90),
	.w8(32'hbbea54fe),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8da585),
	.w1(32'h3b4dc838),
	.w2(32'h3a529b51),
	.w3(32'hba8773ce),
	.w4(32'hb9ece0a7),
	.w5(32'hb9f77a8b),
	.w6(32'hba034dea),
	.w7(32'hbae4454c),
	.w8(32'hb90e9375),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba14bd95),
	.w1(32'hbb2cb9f4),
	.w2(32'hb7cb1e99),
	.w3(32'h3a5e6398),
	.w4(32'h3ac32cc9),
	.w5(32'hba75b4ff),
	.w6(32'hbbb7e95a),
	.w7(32'h398ca5e8),
	.w8(32'hbab558a2),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca1d0de),
	.w1(32'hbc179b60),
	.w2(32'hbb9cdc59),
	.w3(32'hbaed6789),
	.w4(32'h3b865b18),
	.w5(32'h3ba41643),
	.w6(32'hbad2cf64),
	.w7(32'hba012a62),
	.w8(32'hbb9a7073),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbade2f3d),
	.w1(32'h3b0a2604),
	.w2(32'hbae3cb35),
	.w3(32'h39d4242b),
	.w4(32'h3adbd42a),
	.w5(32'h3b0c0147),
	.w6(32'hbc16eaed),
	.w7(32'hbaceeef6),
	.w8(32'h3b8ffdec),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a05e537),
	.w1(32'h3ab06bce),
	.w2(32'hbb229ad5),
	.w3(32'hba0c70b4),
	.w4(32'hbb8fa9fa),
	.w5(32'hbbc3e463),
	.w6(32'hba7d0d84),
	.w7(32'h3a16ff81),
	.w8(32'hb8c2304f),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfc203f),
	.w1(32'hb9a7a4cd),
	.w2(32'h3a82e286),
	.w3(32'h3b566238),
	.w4(32'hbb930ea7),
	.w5(32'hbb1a6b18),
	.w6(32'hbb048bdb),
	.w7(32'h3b15654b),
	.w8(32'h3b3a8d73),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb839fc3),
	.w1(32'hbb50bf68),
	.w2(32'hbb48e6c4),
	.w3(32'hb8cd8d5a),
	.w4(32'h3a31f1f0),
	.w5(32'hbb46f361),
	.w6(32'hbc4a4dcd),
	.w7(32'h3bc763ae),
	.w8(32'h3bffb673),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c811d5e),
	.w1(32'h3b287db1),
	.w2(32'hbaef13e7),
	.w3(32'hbcf1d473),
	.w4(32'hbb0c5878),
	.w5(32'hbb341021),
	.w6(32'hba9b333e),
	.w7(32'hbb824982),
	.w8(32'hbb959692),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d05c244),
	.w1(32'hbc13e22f),
	.w2(32'hbb31014a),
	.w3(32'hbc0b7f86),
	.w4(32'hbbd637b8),
	.w5(32'h3c4864a6),
	.w6(32'hbb5de7d4),
	.w7(32'h3bfb92a0),
	.w8(32'h3b28313c),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3d7413),
	.w1(32'hbb574821),
	.w2(32'h3bda2261),
	.w3(32'h3c452398),
	.w4(32'hb917c94f),
	.w5(32'hbb8dec39),
	.w6(32'hbb9b2a13),
	.w7(32'hbc0174b8),
	.w8(32'hbaecff1b),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b24b00f),
	.w1(32'hbb7cebef),
	.w2(32'hbb716e86),
	.w3(32'h3b94ae3c),
	.w4(32'hb96e35e2),
	.w5(32'h3c29032f),
	.w6(32'hbba65da1),
	.w7(32'h3ba311e5),
	.w8(32'hbc0d2769),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd26cad),
	.w1(32'hbc1aa12b),
	.w2(32'hbb2c1176),
	.w3(32'h3d088033),
	.w4(32'hbc231e09),
	.w5(32'hbb01d21a),
	.w6(32'h3c88c1d9),
	.w7(32'hbbdc9c74),
	.w8(32'h3c849a96),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b30ab7e),
	.w1(32'h3b73ef9f),
	.w2(32'h3ccbb1cd),
	.w3(32'h3c3af744),
	.w4(32'hbbb79518),
	.w5(32'hbbd69461),
	.w6(32'h3b89e1d5),
	.w7(32'h3a1cbb54),
	.w8(32'h3baf0c73),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbacad04),
	.w1(32'hbb80e63a),
	.w2(32'h3b1efced),
	.w3(32'hba10a60a),
	.w4(32'hbb986f9c),
	.w5(32'h3a119f59),
	.w6(32'hba8561ef),
	.w7(32'h3b212a42),
	.w8(32'hbbc5fb51),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a917d92),
	.w1(32'hbc7d36b0),
	.w2(32'hbc092303),
	.w3(32'h3a2dc884),
	.w4(32'h3c02902f),
	.w5(32'hbc258523),
	.w6(32'h3ccf0193),
	.w7(32'h3c9ec3c2),
	.w8(32'hbb7ba625),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3cfc82),
	.w1(32'hbb3bb11f),
	.w2(32'hbb811310),
	.w3(32'hbb733169),
	.w4(32'h3c428cc4),
	.w5(32'hbb8bd4d7),
	.w6(32'h396d988d),
	.w7(32'h3acb70e3),
	.w8(32'hb9c64d08),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae5d9ef),
	.w1(32'h3b5d793d),
	.w2(32'hb857ad7d),
	.w3(32'h3b9f1604),
	.w4(32'h3baa422b),
	.w5(32'hbb803864),
	.w6(32'h3bc6bdca),
	.w7(32'hbc522464),
	.w8(32'h3b7b8803),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d03480d),
	.w1(32'h3bfcf920),
	.w2(32'hbba228b3),
	.w3(32'h3905fbfa),
	.w4(32'hbba8a8eb),
	.w5(32'h3bab8d75),
	.w6(32'hbc17cc23),
	.w7(32'hbc2ac889),
	.w8(32'hbc98e8d6),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba511eb),
	.w1(32'hbb8110f0),
	.w2(32'h3b09d9e4),
	.w3(32'h3a648229),
	.w4(32'hbbb23fbe),
	.w5(32'h3bca70ea),
	.w6(32'hbc227e66),
	.w7(32'hbc0219c5),
	.w8(32'hbbc0322b),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb948d03),
	.w1(32'h34cc3c33),
	.w2(32'h3b576c90),
	.w3(32'hbac33a0f),
	.w4(32'hbc1fda66),
	.w5(32'hbaadc94f),
	.w6(32'hbb37f643),
	.w7(32'h393f373c),
	.w8(32'hbc1b7762),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4147b2),
	.w1(32'hbac4acfb),
	.w2(32'hbba65313),
	.w3(32'hbb590f51),
	.w4(32'hbb5790ac),
	.w5(32'hba6a03e5),
	.w6(32'hbb762866),
	.w7(32'h3b256051),
	.w8(32'hbc603ac0),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc83a108),
	.w1(32'hbbd48ad4),
	.w2(32'hbb9cb92f),
	.w3(32'hbb809b37),
	.w4(32'h3c2868f3),
	.w5(32'hbba20073),
	.w6(32'h3c4ff4f8),
	.w7(32'hbb7a63dd),
	.w8(32'hbaa38058),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb6e6f0),
	.w1(32'hbb912cca),
	.w2(32'h39abf9dd),
	.w3(32'hbba7e079),
	.w4(32'hbb6ba86d),
	.w5(32'hbbf13fc4),
	.w6(32'h3b13adef),
	.w7(32'h3c1f9f70),
	.w8(32'h3afc5c4d),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac8d05f),
	.w1(32'h3b9f5748),
	.w2(32'h3d53280f),
	.w3(32'hbb7188b4),
	.w4(32'h3c0de410),
	.w5(32'h3c3bb5a3),
	.w6(32'hbaedd874),
	.w7(32'h3b03e662),
	.w8(32'hba8b0b8f),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5c51e4),
	.w1(32'h3915196c),
	.w2(32'hbbb752c6),
	.w3(32'h3c59aafe),
	.w4(32'hbbd8eba7),
	.w5(32'hbc352bd3),
	.w6(32'hb8964128),
	.w7(32'hbc478077),
	.w8(32'hbc19a406),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaab607),
	.w1(32'h3d3c9541),
	.w2(32'hbb3744d4),
	.w3(32'hbcda6bba),
	.w4(32'h3c81935b),
	.w5(32'hbbd6743a),
	.w6(32'h3bbe91df),
	.w7(32'hba579881),
	.w8(32'h38405e40),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb5eb0e),
	.w1(32'hbc3f746d),
	.w2(32'hbbd2e5ee),
	.w3(32'hbc7f713f),
	.w4(32'h3a53082f),
	.w5(32'h3a502963),
	.w6(32'hbb81c501),
	.w7(32'hbbf4a042),
	.w8(32'hbbc373e1),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb50f664),
	.w1(32'hbb9524c9),
	.w2(32'hb902e187),
	.w3(32'hbbc26567),
	.w4(32'h3c5bc574),
	.w5(32'h3a32c3ff),
	.w6(32'hb9c004a5),
	.w7(32'hba920655),
	.w8(32'hba6a111f),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf28c1c),
	.w1(32'hbabe98e4),
	.w2(32'h3a0044cf),
	.w3(32'hba6e81ad),
	.w4(32'h3bb473c5),
	.w5(32'h3cd78c9f),
	.w6(32'hbbf5608b),
	.w7(32'hbb59f382),
	.w8(32'hbad15856),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad43e32),
	.w1(32'hb8b2152c),
	.w2(32'h3ae167bd),
	.w3(32'h3b621f24),
	.w4(32'h3afcf010),
	.w5(32'h3acc78f1),
	.w6(32'hba155e16),
	.w7(32'hb8d51501),
	.w8(32'hb7a3a6c3),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b19bda9),
	.w1(32'hbb02f605),
	.w2(32'hbbb3f65e),
	.w3(32'h391cb29c),
	.w4(32'h3df977c7),
	.w5(32'h3c9e4216),
	.w6(32'h3a761a41),
	.w7(32'hbcdcd9f5),
	.w8(32'h3a205d67),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b1e43),
	.w1(32'h3c202f19),
	.w2(32'hbbea512b),
	.w3(32'h3b634c3f),
	.w4(32'hbc3d85c6),
	.w5(32'hbc3d5934),
	.w6(32'hbbbcc835),
	.w7(32'hbc45ff41),
	.w8(32'h3b16f0b8),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba780425),
	.w1(32'hbc794927),
	.w2(32'h3d10e77c),
	.w3(32'hba6f11a2),
	.w4(32'h3a8f96fc),
	.w5(32'hbb143b47),
	.w6(32'hbc414da3),
	.w7(32'h3a3336db),
	.w8(32'h3b5030cf),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbabd273),
	.w1(32'hbc032da3),
	.w2(32'h3bd76ffc),
	.w3(32'h3ab8e47d),
	.w4(32'hbc55b8e8),
	.w5(32'hba2082cd),
	.w6(32'hbc864b66),
	.w7(32'hba6d0c0a),
	.w8(32'hb9000af9),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a56abef),
	.w1(32'hba80f2b1),
	.w2(32'hba2376b0),
	.w3(32'h3b8cfcf9),
	.w4(32'h3afa5da3),
	.w5(32'hbad63a0e),
	.w6(32'hb88af205),
	.w7(32'hba9ce23a),
	.w8(32'hbb245bf9),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb23f20c),
	.w1(32'h3c512bc8),
	.w2(32'hbaabe530),
	.w3(32'h38a93320),
	.w4(32'hbb5617b1),
	.w5(32'hb92c9897),
	.w6(32'h3b08105d),
	.w7(32'hbd26c85c),
	.w8(32'h3a05de45),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b63e32),
	.w1(32'h3860fc07),
	.w2(32'h3aec0d8f),
	.w3(32'h3bb2fc76),
	.w4(32'h3d057772),
	.w5(32'h3afbc6b8),
	.w6(32'h39c381d5),
	.w7(32'h3ad754eb),
	.w8(32'hb9b0cb7c),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ab2c29),
	.w1(32'h3b025abd),
	.w2(32'hbab95682),
	.w3(32'hbb08c66a),
	.w4(32'hbac07034),
	.w5(32'h3b332acf),
	.w6(32'h3d11ac60),
	.w7(32'h3b9828ab),
	.w8(32'hbaf4d680),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d8a8a5),
	.w1(32'h3a20b3a7),
	.w2(32'h3ca76a92),
	.w3(32'h3ac4881b),
	.w4(32'h38a29785),
	.w5(32'hb94ab617),
	.w6(32'hb7efad3e),
	.w7(32'hbad58dee),
	.w8(32'hba886905),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8328541),
	.w1(32'h3b8a9a99),
	.w2(32'hbafa1d6e),
	.w3(32'hbad91970),
	.w4(32'hbaad315c),
	.w5(32'h3aa27a61),
	.w6(32'hb732f7db),
	.w7(32'h3c061d3f),
	.w8(32'hba45e4f6),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba637baf),
	.w1(32'hbb7aa7c2),
	.w2(32'h393a7a5b),
	.w3(32'h3b717c25),
	.w4(32'h3b76f79e),
	.w5(32'hbb9e1cea),
	.w6(32'h3ae609ac),
	.w7(32'h3b236470),
	.w8(32'hba8cc455),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0adcc0),
	.w1(32'hbb2338a4),
	.w2(32'h3b295087),
	.w3(32'h3b0520f3),
	.w4(32'h3b639130),
	.w5(32'h3a18669e),
	.w6(32'h3ad12298),
	.w7(32'hbb807182),
	.w8(32'h3a9b642d),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5d0244),
	.w1(32'h3a2ab8db),
	.w2(32'h39965ba7),
	.w3(32'hba2ad815),
	.w4(32'h3a7f94fd),
	.w5(32'h39e082c5),
	.w6(32'h38875b96),
	.w7(32'h3bfa26a4),
	.w8(32'hb9c7a7ff),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc79494b),
	.w1(32'hb9bc222a),
	.w2(32'h3a7b1f9c),
	.w3(32'hbc4f034c),
	.w4(32'hbb2b8b1b),
	.w5(32'hbb862f13),
	.w6(32'h3b3774ad),
	.w7(32'h3aab2abc),
	.w8(32'h3bb305d8),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fe80b9),
	.w1(32'h3b31fb34),
	.w2(32'h3b7ba464),
	.w3(32'h3b0f68c7),
	.w4(32'hbb5fe2d3),
	.w5(32'hba8a27d0),
	.w6(32'h3c2d1434),
	.w7(32'hbcf31014),
	.w8(32'h3a405481),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0d998e),
	.w1(32'h3aea85e1),
	.w2(32'h3bd5db75),
	.w3(32'h37ae3063),
	.w4(32'h3ba9dce2),
	.w5(32'h3c80382c),
	.w6(32'h3b5feba9),
	.w7(32'hb90a902d),
	.w8(32'hbb6c8fb3),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b278796),
	.w1(32'hba146e0f),
	.w2(32'hbc509b96),
	.w3(32'hbabadc32),
	.w4(32'hbacc4bb7),
	.w5(32'hbaf47747),
	.w6(32'hbb1990a1),
	.w7(32'hb9c9b350),
	.w8(32'hba965b68),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d2a405a),
	.w1(32'h3a97da8a),
	.w2(32'hb8f9a782),
	.w3(32'h3a80f281),
	.w4(32'h3a9c8725),
	.w5(32'hb8c223c5),
	.w6(32'h3cd1a873),
	.w7(32'h3aa80a7c),
	.w8(32'hbb237b7b),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3935284b),
	.w1(32'h3a43908d),
	.w2(32'hba8ee1ee),
	.w3(32'h3a0f1c7f),
	.w4(32'hb92f99e7),
	.w5(32'h3b834eea),
	.w6(32'h3b8c2850),
	.w7(32'hbb201ab8),
	.w8(32'hbbca10c7),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93f1a53),
	.w1(32'h3a917c56),
	.w2(32'h3a9df3d0),
	.w3(32'h399b3f02),
	.w4(32'h3bdb4e9a),
	.w5(32'hbcfd9950),
	.w6(32'hbd31ead7),
	.w7(32'hb92cac97),
	.w8(32'h3bc6afed),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aee44ce),
	.w1(32'h3a805241),
	.w2(32'hbab5189e),
	.w3(32'h3a300c37),
	.w4(32'hba6709a7),
	.w5(32'h3b2e93ad),
	.w6(32'h38c128b6),
	.w7(32'h3b16ff94),
	.w8(32'hb9bfd4c6),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h393b1a09),
	.w1(32'hbc1edd43),
	.w2(32'h370f3149),
	.w3(32'hba0219b6),
	.w4(32'h3b01ec0e),
	.w5(32'hbadea17d),
	.w6(32'hbb16aa6e),
	.w7(32'hbab37fa7),
	.w8(32'h3a58279c),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3c7952),
	.w1(32'h3b88c47e),
	.w2(32'h38a56f67),
	.w3(32'hbcfe040d),
	.w4(32'hbac9b1f6),
	.w5(32'hba6d197a),
	.w6(32'hbae0670c),
	.w7(32'hbd171d3f),
	.w8(32'h3aee1d12),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c93a148),
	.w1(32'hbb448045),
	.w2(32'h3920ba74),
	.w3(32'h398a54af),
	.w4(32'hbb25c59d),
	.w5(32'hbb8309a4),
	.w6(32'h3aae6c49),
	.w7(32'h3d072b07),
	.w8(32'h3c582323),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb847dbe2),
	.w1(32'hbb0d71bc),
	.w2(32'hb9cd5f3a),
	.w3(32'hb9fadbbd),
	.w4(32'hbafd12d7),
	.w5(32'hbb1af1b4),
	.w6(32'hbbaf1d8e),
	.w7(32'h3ca76150),
	.w8(32'h3afa2043),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbe4c9a),
	.w1(32'hbaa8bb30),
	.w2(32'h3a532cc5),
	.w3(32'hb9f7f037),
	.w4(32'hbb8e806d),
	.w5(32'h3adc0630),
	.w6(32'h3cca0a04),
	.w7(32'h3adae547),
	.w8(32'hba46e420),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b105784),
	.w1(32'h392de471),
	.w2(32'h3b154e26),
	.w3(32'h3b811566),
	.w4(32'hbb076982),
	.w5(32'hb92a67d3),
	.w6(32'hb961b4c8),
	.w7(32'h39b04bf6),
	.w8(32'hbb2f58a1),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacf01bb),
	.w1(32'hb8eefb7c),
	.w2(32'hb7e30096),
	.w3(32'hbab862ce),
	.w4(32'h3aa420ce),
	.w5(32'h39aad8f2),
	.w6(32'hbaf94a3d),
	.w7(32'hbb3416ec),
	.w8(32'hbac90bfd),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b587b0),
	.w1(32'hba57734c),
	.w2(32'h3a519455),
	.w3(32'hbb177538),
	.w4(32'hba107c9d),
	.w5(32'hba90e81c),
	.w6(32'hbb973a2f),
	.w7(32'hba53899a),
	.w8(32'h3a85cfc6),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb96c50),
	.w1(32'hbaaf10a0),
	.w2(32'hb9da81c6),
	.w3(32'h3b45282d),
	.w4(32'h3ab98135),
	.w5(32'hb8c250eb),
	.w6(32'hbb267df9),
	.w7(32'hbb1f5fca),
	.w8(32'hb98b0b7c),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab3c9fb),
	.w1(32'h3b22a484),
	.w2(32'hbaa6a6a9),
	.w3(32'hbbd1e0d7),
	.w4(32'hba1932ce),
	.w5(32'h3ab6e361),
	.w6(32'h3ac83978),
	.w7(32'h3bad8b13),
	.w8(32'hbb0a2b1b),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb429f6d),
	.w1(32'h3a907c20),
	.w2(32'h3b3248ba),
	.w3(32'hbba283d4),
	.w4(32'hbbbecc44),
	.w5(32'hba9c60a8),
	.w6(32'h3a56b80f),
	.w7(32'h3b54d356),
	.w8(32'h3b08612c),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90eb569),
	.w1(32'hb83fabd3),
	.w2(32'h3a785242),
	.w3(32'hbac9a47a),
	.w4(32'hbb26f1cf),
	.w5(32'h3b5f95ca),
	.w6(32'hbb3e5afd),
	.w7(32'hbb1709a5),
	.w8(32'h3ab16739),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a77fda5),
	.w1(32'h3b042a89),
	.w2(32'hbb92eda8),
	.w3(32'h3a5fd460),
	.w4(32'h3a84d0e1),
	.w5(32'h3b9c19ec),
	.w6(32'h39597cde),
	.w7(32'hbadb1b4e),
	.w8(32'h3c23ff51),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc278be7),
	.w1(32'hbad43642),
	.w2(32'hba8cd430),
	.w3(32'hb89e1c71),
	.w4(32'h3aebb49e),
	.w5(32'hbac2f778),
	.w6(32'h398c213b),
	.w7(32'hbba11ec0),
	.w8(32'h3c463bd2),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaa205a),
	.w1(32'hbb64d02b),
	.w2(32'h3c94bb09),
	.w3(32'hbadbd110),
	.w4(32'h3965133e),
	.w5(32'h3952c094),
	.w6(32'hbabb2c94),
	.w7(32'hbb2bfbff),
	.w8(32'h3b6a80df),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0e8c0a),
	.w1(32'hba501c01),
	.w2(32'hba06e916),
	.w3(32'h3a77e40b),
	.w4(32'h39dbfc0c),
	.w5(32'hba8b5fc0),
	.w6(32'h3a847838),
	.w7(32'h3b660faf),
	.w8(32'hbbf83b6b),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ae04e4),
	.w1(32'h3bd31b0b),
	.w2(32'h3b86870c),
	.w3(32'h3b73b853),
	.w4(32'h3b66b360),
	.w5(32'h3ba6c6ab),
	.w6(32'h3b6d6bcd),
	.w7(32'h3bb02f25),
	.w8(32'hb90a6085),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb75ce34),
	.w1(32'hbaf17763),
	.w2(32'h38c82f1c),
	.w3(32'h3c787cf9),
	.w4(32'h3b1ad917),
	.w5(32'hba775e2b),
	.w6(32'hb8806d90),
	.w7(32'hb9fb4234),
	.w8(32'hbb4d1853),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ae30f6),
	.w1(32'h3b1181a5),
	.w2(32'hbbb08c26),
	.w3(32'h39dffc2c),
	.w4(32'hba5896b8),
	.w5(32'h3b36023d),
	.w6(32'hbb3f5820),
	.w7(32'hbc5f4498),
	.w8(32'h3a84c323),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabf903f),
	.w1(32'hbb24dc6c),
	.w2(32'h3a7249a5),
	.w3(32'h3af051cc),
	.w4(32'hb9ca17e8),
	.w5(32'h3aa32816),
	.w6(32'hba236c19),
	.w7(32'hbb2c50e4),
	.w8(32'hbabbbf40),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb236eee),
	.w1(32'h3b6684f6),
	.w2(32'hbb166a3a),
	.w3(32'hbb55580e),
	.w4(32'h3b44d128),
	.w5(32'hb9601e2f),
	.w6(32'hbbcdf43b),
	.w7(32'hbb8ffbb4),
	.w8(32'h3ade29da),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9824ad7),
	.w1(32'h3b208f75),
	.w2(32'h3ba26304),
	.w3(32'h3ab12867),
	.w4(32'hb9c98bef),
	.w5(32'hbb5ba656),
	.w6(32'hbb1dfdb0),
	.w7(32'hbaa5bd12),
	.w8(32'h3bbc3bcb),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1114a4),
	.w1(32'h3a0a6af9),
	.w2(32'hbb9e7a43),
	.w3(32'hba9a04ba),
	.w4(32'hbab2e55d),
	.w5(32'hba9ddeb3),
	.w6(32'h39d9526e),
	.w7(32'hb75bd60b),
	.w8(32'h3930e4f1),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fd93c4),
	.w1(32'hbad6b03d),
	.w2(32'h39b367ef),
	.w3(32'h3a17c3ac),
	.w4(32'h3acae783),
	.w5(32'hbba38a09),
	.w6(32'hba5001ca),
	.w7(32'hbad9fc58),
	.w8(32'h3a8ab6cd),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa03e7e),
	.w1(32'h3a3ae0b0),
	.w2(32'h3c1d5d9c),
	.w3(32'hbc0d5ff7),
	.w4(32'h3bc05860),
	.w5(32'h38e419ee),
	.w6(32'h3a206c2a),
	.w7(32'h39417b88),
	.w8(32'hba8a0b43),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb38be62),
	.w1(32'hba9e671f),
	.w2(32'h398911e3),
	.w3(32'hbbd21a16),
	.w4(32'h38967e99),
	.w5(32'hbaca9efc),
	.w6(32'h3792c38b),
	.w7(32'h39b3d013),
	.w8(32'hbbcadd30),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaf9a2a),
	.w1(32'h3b84749e),
	.w2(32'hbb986712),
	.w3(32'h3b920a9c),
	.w4(32'hbb853f22),
	.w5(32'h38bf219c),
	.w6(32'hb8cb77db),
	.w7(32'h3778b9fc),
	.w8(32'hbc1518bd),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7a9a78),
	.w1(32'h3b02f209),
	.w2(32'h3a9dba5d),
	.w3(32'hbbafa828),
	.w4(32'hb84be66b),
	.w5(32'hbaac72f9),
	.w6(32'hbc17dc35),
	.w7(32'hbab8dc76),
	.w8(32'hbb3f4db2),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba07254c),
	.w1(32'hbb18f6cd),
	.w2(32'h3ab65d8a),
	.w3(32'h3b407ef6),
	.w4(32'hbad05b19),
	.w5(32'h39f4dc0d),
	.w6(32'h3a71610d),
	.w7(32'hb8003ea1),
	.w8(32'h3b5c0f6e),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8f121d),
	.w1(32'hbb08bfff),
	.w2(32'h37b181ef),
	.w3(32'h3a1b73de),
	.w4(32'h3b226aac),
	.w5(32'hba0c1bba),
	.w6(32'h3bc335b6),
	.w7(32'h3b2d4157),
	.w8(32'h3a0b623c),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5d98ff),
	.w1(32'h3a0b192d),
	.w2(32'h3b31ad9a),
	.w3(32'hb9d9307f),
	.w4(32'h3ae21ef9),
	.w5(32'h3a647740),
	.w6(32'h3a76ad99),
	.w7(32'hbb1133c3),
	.w8(32'h3b6552ab),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baef899),
	.w1(32'h3c80aa95),
	.w2(32'hbb7631d1),
	.w3(32'h3b881197),
	.w4(32'hb88d43c6),
	.w5(32'h3aa043a0),
	.w6(32'h39bc9509),
	.w7(32'hba7e620b),
	.w8(32'h3a16ac76),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6edb42),
	.w1(32'h3a02a05c),
	.w2(32'h3c015e9d),
	.w3(32'hbabe4dbe),
	.w4(32'hbb88443f),
	.w5(32'h3aef52de),
	.w6(32'h3bbf3186),
	.w7(32'h3acca230),
	.w8(32'h3b067826),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc5b1ee),
	.w1(32'h3b29ea43),
	.w2(32'h3b1614f6),
	.w3(32'h3c02170e),
	.w4(32'hbb11d41d),
	.w5(32'hbada83d6),
	.w6(32'hba94b3de),
	.w7(32'hbac98be5),
	.w8(32'h39e27802),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3577b7),
	.w1(32'hbb316329),
	.w2(32'hba8de650),
	.w3(32'h3b03c4bf),
	.w4(32'hbab3f511),
	.w5(32'h39901eb8),
	.w6(32'hba18dccf),
	.w7(32'h3b697ef4),
	.w8(32'hba87bff7),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc14488),
	.w1(32'hbb00e923),
	.w2(32'h39aef1b6),
	.w3(32'hba837819),
	.w4(32'h3a942951),
	.w5(32'h3aa6038c),
	.w6(32'h3872a131),
	.w7(32'hbb411286),
	.w8(32'hba112323),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f87681),
	.w1(32'h3c24269d),
	.w2(32'h3b693723),
	.w3(32'h39d4fb31),
	.w4(32'h3c0240f3),
	.w5(32'h3b2449e0),
	.w6(32'hbb5d82ba),
	.w7(32'hba71f49e),
	.w8(32'hb947d376),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b16943f),
	.w1(32'h3b8d1ff2),
	.w2(32'h3acacae8),
	.w3(32'hb9db597d),
	.w4(32'h3b5c4e92),
	.w5(32'h3b7e98ca),
	.w6(32'hbad16da8),
	.w7(32'h3bc5b1e3),
	.w8(32'h3b199f1c),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ed54b9),
	.w1(32'hba934658),
	.w2(32'h3b6f530c),
	.w3(32'h3c0054c1),
	.w4(32'hba5e3f2b),
	.w5(32'h3b64ffb1),
	.w6(32'hbab5f48e),
	.w7(32'h3ca2caec),
	.w8(32'hbbb7e90d),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3958872c),
	.w1(32'hbb24e1bf),
	.w2(32'h3aeeb5dd),
	.w3(32'h3b5611c4),
	.w4(32'hba005738),
	.w5(32'h3b3a88a7),
	.w6(32'h3953fdfe),
	.w7(32'h3b28d9c5),
	.w8(32'h3b806524),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba80f9d8),
	.w1(32'h3b6cafed),
	.w2(32'hbc0fc35f),
	.w3(32'hba506985),
	.w4(32'hbac73d55),
	.w5(32'h3a19b911),
	.w6(32'hba8f3f53),
	.w7(32'h3acf36ec),
	.w8(32'hbb21a129),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0736e1),
	.w1(32'hbc49acc7),
	.w2(32'hbb071758),
	.w3(32'hbba3aea2),
	.w4(32'h3b8c5c9f),
	.w5(32'h396c0393),
	.w6(32'h3b9fc440),
	.w7(32'h3ba46512),
	.w8(32'hbb679dca),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a604c7c),
	.w1(32'hbac94bff),
	.w2(32'hbaf6ee44),
	.w3(32'hbb7e4594),
	.w4(32'h3bf98033),
	.w5(32'h3b93fbb1),
	.w6(32'h3aac420e),
	.w7(32'hba40a449),
	.w8(32'hbbf584e1),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba1dff4),
	.w1(32'hbb08e23b),
	.w2(32'hb994c2d6),
	.w3(32'h3b50c7ee),
	.w4(32'h3c2a42d0),
	.w5(32'hb9ced1d1),
	.w6(32'h3b00bf7d),
	.w7(32'h3ac914fb),
	.w8(32'h39f03117),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4651a6),
	.w1(32'h3bc5de82),
	.w2(32'hba8b5e50),
	.w3(32'h3b797646),
	.w4(32'h3b187baf),
	.w5(32'hb827ae8f),
	.w6(32'h39218973),
	.w7(32'h3b8afeed),
	.w8(32'hbb8366ee),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba96ae98),
	.w1(32'hb9f2915e),
	.w2(32'h3828c452),
	.w3(32'hbba958c1),
	.w4(32'h3c830dd7),
	.w5(32'h3ba7058e),
	.w6(32'hbb06e44a),
	.w7(32'hbb628efb),
	.w8(32'h3becc441),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba78f86),
	.w1(32'h3afddf01),
	.w2(32'hbb861b2e),
	.w3(32'h3b2ed97f),
	.w4(32'hbbbe8bc8),
	.w5(32'hbbb3cd6f),
	.w6(32'hbc24b543),
	.w7(32'hbba0b488),
	.w8(32'hb9d33842),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0cca98),
	.w1(32'h3c80d37f),
	.w2(32'h3ab40bc1),
	.w3(32'hbb94ef7b),
	.w4(32'h39f2c917),
	.w5(32'hb8efc027),
	.w6(32'hb996d548),
	.w7(32'hbb8e08e6),
	.w8(32'h3acecfd4),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb244b1),
	.w1(32'hbb32dbc0),
	.w2(32'h3bcb4be5),
	.w3(32'hbb375a7d),
	.w4(32'hba9ba26e),
	.w5(32'h3b546937),
	.w6(32'hbb0f0e0d),
	.w7(32'h3d102505),
	.w8(32'hbb71efb2),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c89517f),
	.w1(32'hbb384870),
	.w2(32'h3b59e8dd),
	.w3(32'h3c5a3ed8),
	.w4(32'h3aca56e6),
	.w5(32'hb8cc33d5),
	.w6(32'hbb2d8828),
	.w7(32'hbb953850),
	.w8(32'h3a0708a2),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb70b67),
	.w1(32'h3915259c),
	.w2(32'h3b906788),
	.w3(32'h3b360025),
	.w4(32'hbb9d6f39),
	.w5(32'hbc24e92f),
	.w6(32'hbb999e4b),
	.w7(32'hb95280a7),
	.w8(32'h3b8bf31e),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cbefc5),
	.w1(32'h3c34d8a6),
	.w2(32'hbc3e1551),
	.w3(32'hbc4948d6),
	.w4(32'h390a9188),
	.w5(32'h3c0f56f7),
	.w6(32'hbaa2605c),
	.w7(32'h3bd16b57),
	.w8(32'h3aa5164b),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2da659),
	.w1(32'h3b188859),
	.w2(32'h3b14e6ba),
	.w3(32'hbafeb979),
	.w4(32'hbb0ebb26),
	.w5(32'hbb0e3aeb),
	.w6(32'hbbb7325a),
	.w7(32'h3cbfb8c3),
	.w8(32'hbc23d7f8),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa31ad1),
	.w1(32'hbb80aa69),
	.w2(32'hb7077666),
	.w3(32'hbb83fc0d),
	.w4(32'hba2456c8),
	.w5(32'hbc25d292),
	.w6(32'hbb6e6143),
	.w7(32'h3b72ec01),
	.w8(32'hb9340bba),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7b3d74),
	.w1(32'hbb08ba0c),
	.w2(32'h3a38cc80),
	.w3(32'h3a951bdd),
	.w4(32'h39f5b532),
	.w5(32'h3b8517df),
	.w6(32'hba822ef9),
	.w7(32'h3a3a5306),
	.w8(32'h3c05e078),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba93b23f),
	.w1(32'hbbb468bf),
	.w2(32'h3c512787),
	.w3(32'hbbd0bd18),
	.w4(32'h3b409378),
	.w5(32'h399368f8),
	.w6(32'h3b128da1),
	.w7(32'h3c09de07),
	.w8(32'h3b8b7ce1),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac65cb7),
	.w1(32'hb9eecfc4),
	.w2(32'hbc28de00),
	.w3(32'h3a8e80c7),
	.w4(32'hbac8ed89),
	.w5(32'hbbb3176e),
	.w6(32'h3b1c5c62),
	.w7(32'h3b452d27),
	.w8(32'h3a9a8e4c),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0a855a),
	.w1(32'h3bd59f37),
	.w2(32'hbb44bc10),
	.w3(32'hbafe37da),
	.w4(32'h3b0762b4),
	.w5(32'hbbb2730e),
	.w6(32'hbbeb18d5),
	.w7(32'h3a9b20ff),
	.w8(32'h3bbcb9e4),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb558536),
	.w1(32'hbb315498),
	.w2(32'h3b77cc31),
	.w3(32'hbbb15445),
	.w4(32'hbb00d81f),
	.w5(32'hba200dc4),
	.w6(32'h3b3be55a),
	.w7(32'hb8a9f39a),
	.w8(32'h3baddce8),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb60dda9),
	.w1(32'h3b2ffbfa),
	.w2(32'hbd446a39),
	.w3(32'hbb5d4374),
	.w4(32'hb90c8fde),
	.w5(32'hbbadb673),
	.w6(32'hbc3c0ea4),
	.w7(32'h381afe68),
	.w8(32'hba40e512),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9840b0),
	.w1(32'hbc034712),
	.w2(32'h3bc6a4d2),
	.w3(32'h3919415c),
	.w4(32'hbc9e54d8),
	.w5(32'hbc02474b),
	.w6(32'hbb5cf506),
	.w7(32'h3b687a74),
	.w8(32'hbaf0ae66),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c03043f),
	.w1(32'h3a29cd1d),
	.w2(32'h3bb01d36),
	.w3(32'hbc80c4e0),
	.w4(32'h3b379f8a),
	.w5(32'hbb04cc8e),
	.w6(32'hbba962f0),
	.w7(32'h3cad749d),
	.w8(32'h3b18cd14),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1f8c7d),
	.w1(32'hbc31d170),
	.w2(32'h3b9af904),
	.w3(32'h3b327e39),
	.w4(32'hbb4274bc),
	.w5(32'h3ca3b377),
	.w6(32'h3988846d),
	.w7(32'h39be3d3b),
	.w8(32'h3bf1a5df),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa7e101),
	.w1(32'hbb4c427c),
	.w2(32'hb91b951b),
	.w3(32'hbc7b309c),
	.w4(32'h3b847508),
	.w5(32'hba2cac17),
	.w6(32'h39ae9a25),
	.w7(32'hbb9ff59f),
	.w8(32'hba0b8f94),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4e8fb0),
	.w1(32'hba88e4d4),
	.w2(32'hbb92bcaf),
	.w3(32'h3aa7cc46),
	.w4(32'h3a14bf7f),
	.w5(32'hbd152e4c),
	.w6(32'hbc01916d),
	.w7(32'h3b3e8067),
	.w8(32'h3c04637d),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c14512f),
	.w1(32'h3afee90c),
	.w2(32'hba840307),
	.w3(32'hbad15cb9),
	.w4(32'h3bc633af),
	.w5(32'hbbc107ff),
	.w6(32'hbbc74e2b),
	.w7(32'hb9890aba),
	.w8(32'h3b12851e),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b83b207),
	.w1(32'h3a931acf),
	.w2(32'hb996eacc),
	.w3(32'h3bc1dad9),
	.w4(32'hbaeff1c9),
	.w5(32'hbb39a7f6),
	.w6(32'hbc196e8e),
	.w7(32'hbaeb3f49),
	.w8(32'h3a5ad924),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1b21f3),
	.w1(32'h3bd9a309),
	.w2(32'hbb49fda6),
	.w3(32'hbc058d88),
	.w4(32'hbb657e85),
	.w5(32'h3a1943ae),
	.w6(32'h3a8318c6),
	.w7(32'h3c538dee),
	.w8(32'hbb2c45f2),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d3312),
	.w1(32'h3b913b98),
	.w2(32'hb94beae9),
	.w3(32'h3b2a6b2c),
	.w4(32'h3b47dadb),
	.w5(32'h3c261d3a),
	.w6(32'hbb873ccc),
	.w7(32'h3a087376),
	.w8(32'h3a251ae4),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae2592c),
	.w1(32'h3b686e11),
	.w2(32'hbbd73ff2),
	.w3(32'h3c058d8e),
	.w4(32'h3cb19b02),
	.w5(32'hbb8951f4),
	.w6(32'hbb2f4629),
	.w7(32'h3b5ce85d),
	.w8(32'hb9b8a6d8),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c52b324),
	.w1(32'h3a37c093),
	.w2(32'hba14c342),
	.w3(32'hbb26d5d7),
	.w4(32'h3a06a4e0),
	.w5(32'h3b791b50),
	.w6(32'h3d2ca9ba),
	.w7(32'hbbbd5233),
	.w8(32'hba50c335),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb995038),
	.w1(32'hbadc8372),
	.w2(32'h3c2174ed),
	.w3(32'h3bc5cc0a),
	.w4(32'hbb3577e4),
	.w5(32'h3b5eca27),
	.w6(32'h3b976c78),
	.w7(32'h3a92f009),
	.w8(32'h3b8b9833),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c34ea30),
	.w1(32'h3a8bfc8b),
	.w2(32'h3c23e14a),
	.w3(32'h3b81ebdb),
	.w4(32'h3b1094ee),
	.w5(32'h3c01818b),
	.w6(32'hbaa8774b),
	.w7(32'hbb1d0c56),
	.w8(32'h3b47e304),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3f5747),
	.w1(32'hbb1fd9ed),
	.w2(32'hbbcdf118),
	.w3(32'h3b07195e),
	.w4(32'hbb3e681b),
	.w5(32'hbae59242),
	.w6(32'h3c45ab37),
	.w7(32'hbb2d3d96),
	.w8(32'hbbddb6b8),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc00e259),
	.w1(32'hbb22cfca),
	.w2(32'h3ae95e32),
	.w3(32'hbb66e4a6),
	.w4(32'h3a092be6),
	.w5(32'hbb28320d),
	.w6(32'hbb13120d),
	.w7(32'h3bbfda62),
	.w8(32'h3bfe3c3c),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb63cdf20),
	.w1(32'h3c2faf27),
	.w2(32'h3ba60b9f),
	.w3(32'h3be82c70),
	.w4(32'h3bb7e4a5),
	.w5(32'hbc0fa090),
	.w6(32'hbb0d446e),
	.w7(32'h3add8922),
	.w8(32'h3c5f48b2),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaf46aa),
	.w1(32'hbb75e690),
	.w2(32'hbb12acf3),
	.w3(32'h3ada6784),
	.w4(32'hbc09da35),
	.w5(32'h3bbdb5d1),
	.w6(32'h3b578c28),
	.w7(32'hba9f0ac3),
	.w8(32'hbae926a8),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba2be65),
	.w1(32'h398eeca5),
	.w2(32'hba8726e7),
	.w3(32'h3ba74552),
	.w4(32'hb99a2612),
	.w5(32'h3c1277e0),
	.w6(32'hba87b728),
	.w7(32'h3cdc6c29),
	.w8(32'h3c21cd01),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc34870f),
	.w1(32'hbaf17e30),
	.w2(32'hbb731bb1),
	.w3(32'h3b84671d),
	.w4(32'hbbcae65b),
	.w5(32'hbb70c86d),
	.w6(32'hbc5b18ed),
	.w7(32'hbab16211),
	.w8(32'h3c02c4b1),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf07349),
	.w1(32'h3af4ad1e),
	.w2(32'h3bbb394c),
	.w3(32'hba018ae2),
	.w4(32'hb7ef848a),
	.w5(32'hbaee792a),
	.w6(32'hbbd867f3),
	.w7(32'h3c70a88a),
	.w8(32'hb88881c1),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb18c2d8),
	.w1(32'hbb882769),
	.w2(32'h3abff628),
	.w3(32'h3a8c5764),
	.w4(32'hbbe16e58),
	.w5(32'hbb54ae0c),
	.w6(32'hb9bcf65e),
	.w7(32'hbb87dc24),
	.w8(32'hba24c9f9),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b21d17c),
	.w1(32'h3a9e99bf),
	.w2(32'hbb522cd5),
	.w3(32'h3a99d1b2),
	.w4(32'h3b420c87),
	.w5(32'h399de493),
	.w6(32'hb919d701),
	.w7(32'h39cc9ca7),
	.w8(32'h3b6390b3),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6978c0),
	.w1(32'h3941457a),
	.w2(32'hbb93802a),
	.w3(32'h39371b19),
	.w4(32'hbb6ffc9d),
	.w5(32'h3c218a62),
	.w6(32'h3bfea1ff),
	.w7(32'h3b5eed59),
	.w8(32'h3b7b3a61),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad624a6),
	.w1(32'hbbbd2f42),
	.w2(32'h3b8b0370),
	.w3(32'hbbccf00e),
	.w4(32'hba13fd30),
	.w5(32'hbbab9e14),
	.w6(32'hbb00150c),
	.w7(32'hbc14811a),
	.w8(32'h3c69d083),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c817bda),
	.w1(32'h3923d8d8),
	.w2(32'h3aaca5a5),
	.w3(32'h3a7b27f6),
	.w4(32'h3bebad50),
	.w5(32'h3bb5287e),
	.w6(32'h3ad8adfc),
	.w7(32'hbb823869),
	.w8(32'h3b702881),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae2f997),
	.w1(32'hbab12674),
	.w2(32'hbbba4af6),
	.w3(32'h3862ddaa),
	.w4(32'hbb0de3e6),
	.w5(32'h3b97b7a7),
	.w6(32'hbba7f737),
	.w7(32'hbb2d3cc2),
	.w8(32'h3a6706d7),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaec450d),
	.w1(32'h3aa75b19),
	.w2(32'h3ba719bf),
	.w3(32'hba666535),
	.w4(32'hbba76a88),
	.w5(32'h3b2298f6),
	.w6(32'hbb4d646c),
	.w7(32'h3b9f240a),
	.w8(32'hb953eed6),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36c2fd9d),
	.w1(32'h39a42dc1),
	.w2(32'h3b7772f4),
	.w3(32'h3bc6810b),
	.w4(32'h3a2388a1),
	.w5(32'hbc0857b3),
	.w6(32'h3af8b395),
	.w7(32'hba242d84),
	.w8(32'h3bc57839),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb731d55),
	.w1(32'hba5c9494),
	.w2(32'h3a2adf46),
	.w3(32'h3c2d6151),
	.w4(32'h3aea6ace),
	.w5(32'h3a8e3bd3),
	.w6(32'hbbfb4178),
	.w7(32'h3c12e309),
	.w8(32'hbbdce0e6),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7b8a48),
	.w1(32'hbb859e4b),
	.w2(32'hba07d312),
	.w3(32'h3be7ce23),
	.w4(32'h3bb4f695),
	.w5(32'hba8b2904),
	.w6(32'hbc28457b),
	.w7(32'hbac1c69e),
	.w8(32'h3bae4877),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c17e9c0),
	.w1(32'h3a149428),
	.w2(32'hb9ea91c0),
	.w3(32'h3b4af9f3),
	.w4(32'h3a91b12f),
	.w5(32'hbb69cc04),
	.w6(32'h3c2d52b3),
	.w7(32'hbb7a61dc),
	.w8(32'hbb8d3f16),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb676c98),
	.w1(32'h3c926d41),
	.w2(32'hbabde6b0),
	.w3(32'h3aebd94f),
	.w4(32'hbae02612),
	.w5(32'hbb8572ca),
	.w6(32'h3c0a08f9),
	.w7(32'hbb090305),
	.w8(32'h3b77130b),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdfc699),
	.w1(32'hbb8f759f),
	.w2(32'hbb74f1df),
	.w3(32'h3978fe56),
	.w4(32'h3baf8a26),
	.w5(32'h3c6ee9fc),
	.w6(32'hbb1ee03c),
	.w7(32'hbb947592),
	.w8(32'h3942a8d9),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b04025),
	.w1(32'hbc5475e3),
	.w2(32'hbb3e3da9),
	.w3(32'h3b8dac9b),
	.w4(32'h3bf9d931),
	.w5(32'h3af6a799),
	.w6(32'hbbdba879),
	.w7(32'h3c3c00be),
	.w8(32'hb78f8f00),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b345646),
	.w1(32'hbc112747),
	.w2(32'h3a05b81a),
	.w3(32'h3c1964e8),
	.w4(32'h3a8171a3),
	.w5(32'hbbad1eb5),
	.w6(32'h3c2a8fae),
	.w7(32'h3b42bcb0),
	.w8(32'hbb51ea93),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b761aad),
	.w1(32'hbbbfe972),
	.w2(32'h3b6b8157),
	.w3(32'hb5a61792),
	.w4(32'hbb9bf447),
	.w5(32'h3bb040ed),
	.w6(32'h3b416953),
	.w7(32'hbc3863ac),
	.w8(32'hbadd151f),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6f0f09),
	.w1(32'hba940d4f),
	.w2(32'h3b688da4),
	.w3(32'h3cb9b9e2),
	.w4(32'hbb2c7ca2),
	.w5(32'h3bbf38b1),
	.w6(32'h3b87ba64),
	.w7(32'hbabdc7cb),
	.w8(32'hbaadbe45),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2e4883),
	.w1(32'hb9286710),
	.w2(32'hbb1ac621),
	.w3(32'h3aeb37aa),
	.w4(32'h3c4891ba),
	.w5(32'hbb63fbd6),
	.w6(32'h3bc9ca7d),
	.w7(32'h3c07592c),
	.w8(32'h3b4a0e4f),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c119cfb),
	.w1(32'h3c2d33f6),
	.w2(32'h3c99c8b7),
	.w3(32'hb9fcaa3d),
	.w4(32'h3a3e1867),
	.w5(32'hbb7782bd),
	.w6(32'hbb0f4ff1),
	.w7(32'hbc042226),
	.w8(32'hbbc0c82e),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule