module layer_8_featuremap_10(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc717290),
	.w1(32'hbb0fbc90),
	.w2(32'hbb953edd),
	.w3(32'h3c9ecc78),
	.w4(32'hbb2ff88d),
	.w5(32'hbb816be3),
	.w6(32'h3c88798a),
	.w7(32'hb9b4a500),
	.w8(32'hbb063832),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4113a3),
	.w1(32'hbadcf16c),
	.w2(32'hbb88ed25),
	.w3(32'hbac13136),
	.w4(32'hbb95da51),
	.w5(32'hbbe7bbdb),
	.w6(32'hb986f31b),
	.w7(32'hbbc1fed4),
	.w8(32'hbb2e4420),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb89c7f4),
	.w1(32'hbb80cd1e),
	.w2(32'hbc01af64),
	.w3(32'hbbc488eb),
	.w4(32'hba557625),
	.w5(32'hbb4bcd78),
	.w6(32'hbb690201),
	.w7(32'hba85be67),
	.w8(32'h3ae03512),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5a6155),
	.w1(32'hbad12be7),
	.w2(32'hbc29a4c4),
	.w3(32'hbb831536),
	.w4(32'h3ba1ad4e),
	.w5(32'h3b217624),
	.w6(32'hbaf6cd51),
	.w7(32'hba97c4b3),
	.w8(32'h3ad8dabd),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0a9bc9),
	.w1(32'hb77b6fb0),
	.w2(32'hbb0af985),
	.w3(32'h3b326958),
	.w4(32'h3b205d2a),
	.w5(32'h3a0ee93f),
	.w6(32'h3b9d5b1f),
	.w7(32'h3b5b5aeb),
	.w8(32'h3a8a4c85),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8e3597),
	.w1(32'hba8d6e9d),
	.w2(32'hbabd11c3),
	.w3(32'h3a48853e),
	.w4(32'hbb1a95bc),
	.w5(32'hb9847c76),
	.w6(32'h3a7c27c8),
	.w7(32'hbab535eb),
	.w8(32'hba3eb50d),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabf4cb7),
	.w1(32'hb9228854),
	.w2(32'hb9d7fad3),
	.w3(32'hb9d17a65),
	.w4(32'hb80b86e7),
	.w5(32'hbaa4600f),
	.w6(32'h3ac8219a),
	.w7(32'hb9aca58a),
	.w8(32'hbad9d9f9),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9f19d0),
	.w1(32'hbad5c66f),
	.w2(32'h3a279158),
	.w3(32'hbb0581d2),
	.w4(32'hba8f841e),
	.w5(32'hb7f0635c),
	.w6(32'hbac64de9),
	.w7(32'h3a160677),
	.w8(32'h3b61f714),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba823127),
	.w1(32'hba83aef5),
	.w2(32'h378b087e),
	.w3(32'h3b1ee0cc),
	.w4(32'h3a303700),
	.w5(32'h3ac83543),
	.w6(32'hb9b34a5e),
	.w7(32'hba00f2bd),
	.w8(32'h39b76650),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389cd024),
	.w1(32'h3a3eee88),
	.w2(32'hb800f9af),
	.w3(32'h3a802bbb),
	.w4(32'h3b5347e4),
	.w5(32'h3b3c7b0a),
	.w6(32'h3aecda99),
	.w7(32'hb9ba6ac1),
	.w8(32'h3b195c5c),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2d3e93),
	.w1(32'h3981e65e),
	.w2(32'hba967957),
	.w3(32'h3b78c6d5),
	.w4(32'h3a8ad767),
	.w5(32'h3a34b24c),
	.w6(32'h3b50e597),
	.w7(32'h3a728c1e),
	.w8(32'h3a2bdc1b),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba306647),
	.w1(32'hba4b3bbb),
	.w2(32'hb92abb28),
	.w3(32'h3a531dab),
	.w4(32'hba37548d),
	.w5(32'h3b21016d),
	.w6(32'h3ab293a5),
	.w7(32'hbb48652f),
	.w8(32'hbaa3f53f),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb959fb6d),
	.w1(32'h3afaa20e),
	.w2(32'h3aed77f2),
	.w3(32'h3b81699b),
	.w4(32'hba9692d6),
	.w5(32'hb892458a),
	.w6(32'h3ac36780),
	.w7(32'hb9698124),
	.w8(32'h39b0e4b3),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbace735c),
	.w1(32'hbb13d42e),
	.w2(32'h38e8c52e),
	.w3(32'hba8de9dd),
	.w4(32'hbab31f75),
	.w5(32'h3b001b5e),
	.w6(32'h39c1331d),
	.w7(32'h3a923973),
	.w8(32'h3b901bb7),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af2b45b),
	.w1(32'h39a9c8af),
	.w2(32'hb941c24a),
	.w3(32'h3b938fca),
	.w4(32'h395800a4),
	.w5(32'hb9c3d418),
	.w6(32'h3bced162),
	.w7(32'hb9ad1a56),
	.w8(32'hb9fe8297),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4e0b72),
	.w1(32'h39555236),
	.w2(32'hb9a3b084),
	.w3(32'hbaa8412b),
	.w4(32'hba352374),
	.w5(32'hb91a9a1e),
	.w6(32'hbac1cb04),
	.w7(32'hbac0dfd7),
	.w8(32'h3a8343e1),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba749957),
	.w1(32'hba908ce8),
	.w2(32'h3aad9827),
	.w3(32'hb8ddc069),
	.w4(32'hba9911b3),
	.w5(32'h3ab8367a),
	.w6(32'h3aec8e48),
	.w7(32'hbaa59949),
	.w8(32'hba4d733f),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0ceac3),
	.w1(32'h3884a5be),
	.w2(32'h3a81a618),
	.w3(32'h3b9ed7e3),
	.w4(32'hbab11693),
	.w5(32'h3aa0bba1),
	.w6(32'h3a5fb39d),
	.w7(32'h399db851),
	.w8(32'h3addd8f3),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a496be3),
	.w1(32'h3a00a79d),
	.w2(32'h3a2a33ec),
	.w3(32'h3b1c6583),
	.w4(32'h3ae15d53),
	.w5(32'h3b415e25),
	.w6(32'h3b876165),
	.w7(32'h3a322733),
	.w8(32'h3a858668),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7af12b7),
	.w1(32'h3add2101),
	.w2(32'h3b322634),
	.w3(32'h3a97f121),
	.w4(32'h3b44a765),
	.w5(32'h3b21c81e),
	.w6(32'h3b5df336),
	.w7(32'h3b1628d2),
	.w8(32'h3a4ea19d),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3816ca3f),
	.w1(32'hb940ddd4),
	.w2(32'h3acd9060),
	.w3(32'hb9f26296),
	.w4(32'h39e68021),
	.w5(32'h3b7dd557),
	.w6(32'hb8c94585),
	.w7(32'h3ada43b5),
	.w8(32'h3ba015bc),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9c4298),
	.w1(32'hb89de92d),
	.w2(32'h3b9b579e),
	.w3(32'h3b51fad1),
	.w4(32'hbac2b734),
	.w5(32'h3a32b0a9),
	.w6(32'h3bbb4b36),
	.w7(32'hba88d6ee),
	.w8(32'h38c90105),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3f311c),
	.w1(32'h374689e3),
	.w2(32'hb9931fa2),
	.w3(32'h3b23e44d),
	.w4(32'hba1b720d),
	.w5(32'h3a94d33a),
	.w6(32'h3ae64351),
	.w7(32'h3aca4776),
	.w8(32'hb830dbaf),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbace94b1),
	.w1(32'hba870b4c),
	.w2(32'hba986489),
	.w3(32'hbac47a20),
	.w4(32'hbabb834c),
	.w5(32'hbaeb873f),
	.w6(32'hbaa1484a),
	.w7(32'hba5abd65),
	.w8(32'hbb289fe5),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8e8cba),
	.w1(32'h3b2baba3),
	.w2(32'h3b13ecd0),
	.w3(32'hbb114478),
	.w4(32'h3b004f7a),
	.w5(32'h3bcf6b9d),
	.w6(32'hbb77520b),
	.w7(32'h3b207744),
	.w8(32'h3b9b6f4a),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b69131e),
	.w1(32'h3939c237),
	.w2(32'hbab169a2),
	.w3(32'h3b8f0513),
	.w4(32'h3a278412),
	.w5(32'hb8dec16a),
	.w6(32'h3b182d29),
	.w7(32'hb8f0baed),
	.w8(32'hbb03977d),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba83dd1d),
	.w1(32'h398e4c8c),
	.w2(32'hb98b92b5),
	.w3(32'hbb1f92a7),
	.w4(32'hb9d3ec6b),
	.w5(32'hb8ed7983),
	.w6(32'hbb4d2f08),
	.w7(32'hb954f1d9),
	.w8(32'h39ac3332),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9898b51),
	.w1(32'hbafef3a6),
	.w2(32'hbb3b2153),
	.w3(32'h3b07cd87),
	.w4(32'h39e0ee39),
	.w5(32'hbadb881b),
	.w6(32'h3a825e3f),
	.w7(32'hbacb664f),
	.w8(32'hbb343e3f),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa6b00a),
	.w1(32'h3a079290),
	.w2(32'h3a7beb06),
	.w3(32'hbb5bb00f),
	.w4(32'h3a8d5ca5),
	.w5(32'h3ab9dc77),
	.w6(32'h3953e00f),
	.w7(32'hba57baa3),
	.w8(32'h396dd8bf),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabb69de),
	.w1(32'hba1a5984),
	.w2(32'h3a7bb6fd),
	.w3(32'hba2b6098),
	.w4(32'hba41079c),
	.w5(32'h39f2132e),
	.w6(32'h39de0fa9),
	.w7(32'hb91d0dfc),
	.w8(32'h3aa1724d),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa07ec9),
	.w1(32'hbb55991c),
	.w2(32'hbaed0f03),
	.w3(32'hbab773ed),
	.w4(32'hbba30f65),
	.w5(32'hbb539760),
	.w6(32'hbaa5e960),
	.w7(32'hbb86c82f),
	.w8(32'hbb48b182),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba56768d),
	.w1(32'h37b5c0e4),
	.w2(32'hb9cf3745),
	.w3(32'hbb03c8f2),
	.w4(32'h3798edb9),
	.w5(32'hba3c94f2),
	.w6(32'hbb508a02),
	.w7(32'hbae1fdcd),
	.w8(32'hbb2302b9),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab7957c),
	.w1(32'hb9a3ca8a),
	.w2(32'hb8965c65),
	.w3(32'hbb057760),
	.w4(32'hb93698bb),
	.w5(32'h388a8310),
	.w6(32'hbb2f9107),
	.w7(32'h38797f26),
	.w8(32'h399224f9),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3913886a),
	.w1(32'hbaf2ef8b),
	.w2(32'hbb00fadb),
	.w3(32'h3a03316c),
	.w4(32'hba8b7baa),
	.w5(32'hbabb8605),
	.w6(32'h3a7ba06e),
	.w7(32'hba9b12fe),
	.w8(32'hbae8f4a5),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa7ed78),
	.w1(32'h39dcff67),
	.w2(32'h3b15db1b),
	.w3(32'hb9de8419),
	.w4(32'h3a04b9e4),
	.w5(32'h3b06fab2),
	.w6(32'hb9655c32),
	.w7(32'h39c7df3d),
	.w8(32'h3ad6a610),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7f34c21),
	.w1(32'h39a6d3d2),
	.w2(32'h3aa0f6dd),
	.w3(32'h3a511204),
	.w4(32'hb9e5532b),
	.w5(32'h3a0e3647),
	.w6(32'h3a8cd144),
	.w7(32'hba5820df),
	.w8(32'hb803baf9),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93f5ec1),
	.w1(32'hbaf182ca),
	.w2(32'hbb7297f6),
	.w3(32'hb9109357),
	.w4(32'hbb4f09fe),
	.w5(32'hbbb946b4),
	.w6(32'hbac0fdc3),
	.w7(32'hbb877e7a),
	.w8(32'hbba0cf5d),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3218c2),
	.w1(32'h3b319422),
	.w2(32'h3b5110d9),
	.w3(32'hbb804860),
	.w4(32'h3b384dcf),
	.w5(32'h3b4a64af),
	.w6(32'hbb431e59),
	.w7(32'h3b51dccc),
	.w8(32'h3b494e2a),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad59f28),
	.w1(32'hba3308ca),
	.w2(32'h38d7cf88),
	.w3(32'hba8a92ae),
	.w4(32'hbaf93162),
	.w5(32'h39fea30b),
	.w6(32'hbaea7aff),
	.w7(32'hbaba3a10),
	.w8(32'hba570aed),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb07547c),
	.w1(32'hba2e1df4),
	.w2(32'h39b17f5c),
	.w3(32'hbb173a6d),
	.w4(32'h39b8b9b9),
	.w5(32'hb98ee867),
	.w6(32'hba91d435),
	.w7(32'hba468e5d),
	.w8(32'hba94c4e5),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e43f7b),
	.w1(32'hba86d4cd),
	.w2(32'h399bd52e),
	.w3(32'hba723240),
	.w4(32'h3a8e7431),
	.w5(32'h3b45e084),
	.w6(32'hb93e880e),
	.w7(32'h3ac4d4d2),
	.w8(32'h3b20fd06),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb938b719),
	.w1(32'hba3f6bf3),
	.w2(32'h3a2cd958),
	.w3(32'h3ae1d7f5),
	.w4(32'hb994986c),
	.w5(32'h3ac747ab),
	.w6(32'h3a3c534e),
	.w7(32'h3a4b7dc9),
	.w8(32'h3b150c73),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b117117),
	.w1(32'h3a3dcbb7),
	.w2(32'h3aaf102e),
	.w3(32'h3b552243),
	.w4(32'h3aa19a1f),
	.w5(32'h3ad3fc67),
	.w6(32'h3b829398),
	.w7(32'h39a1f8b7),
	.w8(32'h3993d9e2),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39332d3b),
	.w1(32'hbb592035),
	.w2(32'hbb037570),
	.w3(32'h39fc1dd7),
	.w4(32'hbb9ad4d0),
	.w5(32'hbb36873b),
	.w6(32'h3a0de4de),
	.w7(32'hbb081e37),
	.w8(32'hbb296f4d),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac5ff36),
	.w1(32'h39d1466d),
	.w2(32'h3ac26472),
	.w3(32'hbafa17f8),
	.w4(32'h3b07dd3d),
	.w5(32'h3b491b07),
	.w6(32'hbac1571d),
	.w7(32'h3b424431),
	.w8(32'h3b8273f2),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a776a44),
	.w1(32'h3a8a2a44),
	.w2(32'hba3256ca),
	.w3(32'h3b199e50),
	.w4(32'h3b2db856),
	.w5(32'h3ada01fe),
	.w6(32'h3b8204b7),
	.w7(32'h38573b78),
	.w8(32'h392b244d),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf4c2a0),
	.w1(32'hba36e8f9),
	.w2(32'h3a94bc86),
	.w3(32'hb9d2c1f7),
	.w4(32'hb974d844),
	.w5(32'h3ace2920),
	.w6(32'hb9d2acf8),
	.w7(32'hbb031289),
	.w8(32'h3a2e2386),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397d2893),
	.w1(32'hbae4f176),
	.w2(32'h3921c029),
	.w3(32'h3b4a589b),
	.w4(32'h38adb094),
	.w5(32'h384697ae),
	.w6(32'h3a8a3ee0),
	.w7(32'h3b114627),
	.w8(32'hb8fcc6b5),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39962e4b),
	.w1(32'h3a7ec8fb),
	.w2(32'hb9a3208d),
	.w3(32'hbb093ff7),
	.w4(32'h3a207586),
	.w5(32'hba35382d),
	.w6(32'hba6ddee8),
	.w7(32'h390267e0),
	.w8(32'hba8c43f3),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9ad05c),
	.w1(32'h39eb0376),
	.w2(32'hba4cff01),
	.w3(32'hbb0ab6d5),
	.w4(32'h3aecf46a),
	.w5(32'h3ab743b1),
	.w6(32'hbadc0942),
	.w7(32'hb90e74d5),
	.w8(32'h3a37550d),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb87bb71),
	.w1(32'hbb21cd0e),
	.w2(32'hba90a310),
	.w3(32'hbabdf41e),
	.w4(32'hbaec13ae),
	.w5(32'hba611556),
	.w6(32'hba90f878),
	.w7(32'hbb4e31fb),
	.w8(32'hbab73cc2),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba93ec37),
	.w1(32'h3a950f21),
	.w2(32'h3b5cd054),
	.w3(32'hba2d965b),
	.w4(32'h39ff1a1d),
	.w5(32'h3b47988d),
	.w6(32'h3a8c815b),
	.w7(32'h3b49c313),
	.w8(32'h3ba49f02),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7bca31),
	.w1(32'hbac66505),
	.w2(32'hb963517f),
	.w3(32'h3aa016ac),
	.w4(32'hba400ef2),
	.w5(32'hba37011f),
	.w6(32'h3b14bdb3),
	.w7(32'h3abaad10),
	.w8(32'h3ae44668),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac2f7ab),
	.w1(32'h3b626bb1),
	.w2(32'hba02d7f3),
	.w3(32'h3ae68d28),
	.w4(32'h399aceed),
	.w5(32'h3b04f157),
	.w6(32'hba4e2a07),
	.w7(32'hbab06a83),
	.w8(32'hb975d327),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaed5693),
	.w1(32'hba36741b),
	.w2(32'hbb591ad3),
	.w3(32'h3b38f2c5),
	.w4(32'h3a33bfeb),
	.w5(32'hb9f4e36f),
	.w6(32'h3b22913f),
	.w7(32'h3ad0a978),
	.w8(32'h3b4e3bd1),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcb8a6e),
	.w1(32'hbac65c5f),
	.w2(32'hba846325),
	.w3(32'hbb2fec5c),
	.w4(32'h397360c3),
	.w5(32'h3a978a5a),
	.w6(32'h3abd4eb3),
	.w7(32'hba041097),
	.w8(32'h394a1ddd),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39174112),
	.w1(32'h3984219c),
	.w2(32'hb612df0b),
	.w3(32'h3a32e4fc),
	.w4(32'h3a4141b5),
	.w5(32'h3846fc26),
	.w6(32'h3a624d11),
	.w7(32'h38e25e99),
	.w8(32'h39be4c27),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a4d1dd),
	.w1(32'hbacd2d13),
	.w2(32'hb9a793fb),
	.w3(32'hba90061b),
	.w4(32'hbafb699d),
	.w5(32'hb99ee67a),
	.w6(32'hba08f7f7),
	.w7(32'hbb3137a6),
	.w8(32'hb7b09d69),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba05735f),
	.w1(32'h382c9eed),
	.w2(32'hb9c91841),
	.w3(32'hbab77567),
	.w4(32'h38261a1a),
	.w5(32'h38345c91),
	.w6(32'h3837e8ae),
	.w7(32'hb9f8124e),
	.w8(32'h39800b0c),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba74913e),
	.w1(32'h3ae27714),
	.w2(32'h3ad68a00),
	.w3(32'hb8d5b624),
	.w4(32'h3abb7a87),
	.w5(32'h3b67b550),
	.w6(32'h3a0dbb4e),
	.w7(32'h3a56afa8),
	.w8(32'h3b9e1624),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3afc43),
	.w1(32'h3a9d506b),
	.w2(32'hba3b328f),
	.w3(32'h3b446851),
	.w4(32'hb950f869),
	.w5(32'hbaa29f41),
	.w6(32'h3af51450),
	.w7(32'hbab9130d),
	.w8(32'h3b24e947),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8859f8),
	.w1(32'hbad9bfa8),
	.w2(32'hba37c4c9),
	.w3(32'h3b64617b),
	.w4(32'hbb0902f3),
	.w5(32'hb9cff692),
	.w6(32'h3c347744),
	.w7(32'hbae96087),
	.w8(32'hba9921aa),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1e6513),
	.w1(32'h3aba7442),
	.w2(32'h3a45e696),
	.w3(32'hba51a71d),
	.w4(32'h3afeaa5a),
	.w5(32'h3aed2223),
	.w6(32'hbab86345),
	.w7(32'h3ae3c2d2),
	.w8(32'h3ad71dbb),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a72f371),
	.w1(32'h3acb743f),
	.w2(32'hba8b2c40),
	.w3(32'h3a92f381),
	.w4(32'h3b530dda),
	.w5(32'h3ae093f8),
	.w6(32'h3b0d35d0),
	.w7(32'h3acf7d5f),
	.w8(32'h3b4cade8),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba37dff5),
	.w1(32'h399efb0b),
	.w2(32'hba99b595),
	.w3(32'h3b57d46b),
	.w4(32'hb80e2190),
	.w5(32'hba033135),
	.w6(32'h3b14046f),
	.w7(32'h39babc19),
	.w8(32'h39e11d94),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f3cdb3),
	.w1(32'h3953ed43),
	.w2(32'hb93e81d9),
	.w3(32'h3ad96320),
	.w4(32'h384ea213),
	.w5(32'h3988fa75),
	.w6(32'h3b1b16c4),
	.w7(32'h39e4a234),
	.w8(32'h3a137522),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ada5537),
	.w1(32'h3a217727),
	.w2(32'h3adba235),
	.w3(32'h3b31a1e5),
	.w4(32'h3acaa838),
	.w5(32'h3b824ce2),
	.w6(32'h3b636605),
	.w7(32'h3b1667f8),
	.w8(32'h3b7ec502),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae1f08e),
	.w1(32'h3a6a58fb),
	.w2(32'h3b2c5d36),
	.w3(32'h3b81dbd9),
	.w4(32'h3b0adfd6),
	.w5(32'h3b8db355),
	.w6(32'h3b9dffc2),
	.w7(32'h3b48add7),
	.w8(32'h3bb7dff5),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8899e4),
	.w1(32'hb9ad21ba),
	.w2(32'hbaa6954f),
	.w3(32'h3bb9f18a),
	.w4(32'hbaf53de4),
	.w5(32'hbada96a9),
	.w6(32'h3bd0c46e),
	.w7(32'hba517b1c),
	.w8(32'h37e9867e),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb117234),
	.w1(32'h3a329c18),
	.w2(32'hbb9cda41),
	.w3(32'hb9314112),
	.w4(32'hbbfb580a),
	.w5(32'hba09aade),
	.w6(32'h3a6ab16b),
	.w7(32'hbc02d0fa),
	.w8(32'hbb0ac56b),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2d73a4),
	.w1(32'hba1b8f09),
	.w2(32'h3ac12f83),
	.w3(32'hb9fbda08),
	.w4(32'hbb093bde),
	.w5(32'hbb4a68f2),
	.w6(32'hbc03cace),
	.w7(32'hbbe210fb),
	.w8(32'hbaa2a95c),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaffcab0),
	.w1(32'hbc95d720),
	.w2(32'h3b89cf2e),
	.w3(32'h398670df),
	.w4(32'hbaa9db45),
	.w5(32'hbc0506f3),
	.w6(32'hba70d593),
	.w7(32'h3be8dfc2),
	.w8(32'hbc9cb1ca),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9595008),
	.w1(32'hbb895234),
	.w2(32'hbaeb9f5a),
	.w3(32'h3a638dcd),
	.w4(32'hbb5e4ad9),
	.w5(32'hbae4bf6b),
	.w6(32'hba5c0d07),
	.w7(32'h39e45aa6),
	.w8(32'hb9eee59f),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6c7039),
	.w1(32'hbbd4ed45),
	.w2(32'h3c0b4b86),
	.w3(32'hbb0367a8),
	.w4(32'hbc25eec6),
	.w5(32'h38e359d1),
	.w6(32'hbb44337e),
	.w7(32'h3bdacdea),
	.w8(32'hbc5aab4c),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c586ca1),
	.w1(32'hbb1de9e0),
	.w2(32'h3ab385e1),
	.w3(32'h3b4b06ab),
	.w4(32'hbb267395),
	.w5(32'hbb8b1120),
	.w6(32'h3bee547b),
	.w7(32'h3bbd7b84),
	.w8(32'h3b18f685),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0d9811),
	.w1(32'hbc5576d5),
	.w2(32'h38589585),
	.w3(32'hba7f5db6),
	.w4(32'hbc62772b),
	.w5(32'hbbf355be),
	.w6(32'hba08c789),
	.w7(32'h3c275528),
	.w8(32'hbd027837),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb3333f),
	.w1(32'hbc46a050),
	.w2(32'h3cb62dc3),
	.w3(32'hbc592287),
	.w4(32'hbcd7383a),
	.w5(32'h3cfff2c0),
	.w6(32'hbbe2cbee),
	.w7(32'h3c74cd97),
	.w8(32'hbcd3bccc),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb272b1),
	.w1(32'hbb84ee0c),
	.w2(32'hbb18b1e1),
	.w3(32'h3c2c4967),
	.w4(32'hbb4befa5),
	.w5(32'h3affbdea),
	.w6(32'h3c008569),
	.w7(32'h3ba63e39),
	.w8(32'h3b2c7aad),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1172e8),
	.w1(32'hbae0e194),
	.w2(32'h3af05c13),
	.w3(32'hbb8ab95b),
	.w4(32'h3a683a1f),
	.w5(32'hbb100416),
	.w6(32'h3b90a61b),
	.w7(32'hbb978514),
	.w8(32'hbb353c59),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4d87be),
	.w1(32'hbb3b2dfd),
	.w2(32'hba9e1691),
	.w3(32'h399d0daf),
	.w4(32'h3bdcdd23),
	.w5(32'hb9cfc6fe),
	.w6(32'hbba512f8),
	.w7(32'h3bbd562f),
	.w8(32'h3affb769),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae42b4d),
	.w1(32'hbbd17c31),
	.w2(32'hbc0d7993),
	.w3(32'hbbc6a9bd),
	.w4(32'h3c2edecb),
	.w5(32'hbc23cf75),
	.w6(32'hbb0b9589),
	.w7(32'hbb55130a),
	.w8(32'hbb9bcc6b),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2ccec5),
	.w1(32'h3a48ef27),
	.w2(32'h3b46aa0d),
	.w3(32'h3bf53f42),
	.w4(32'h3ada57d8),
	.w5(32'h3b6f35f3),
	.w6(32'hbc1d7be4),
	.w7(32'h3b88be1b),
	.w8(32'h3a82c02b),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389286d5),
	.w1(32'h3bb03b8a),
	.w2(32'hbd4547ff),
	.w3(32'h3b2689db),
	.w4(32'h3d0e1fb1),
	.w5(32'hbce56881),
	.w6(32'h3bab0cf7),
	.w7(32'hbc798f6a),
	.w8(32'h3d763c4d),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d2268ba),
	.w1(32'hb9b8ab6b),
	.w2(32'h3c01f7f9),
	.w3(32'hbb291e8b),
	.w4(32'h3a2c2308),
	.w5(32'h3b3ca56a),
	.w6(32'hbd718c65),
	.w7(32'hbb2f23a0),
	.w8(32'h39046f29),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b87dcae),
	.w1(32'hbc0ebdd5),
	.w2(32'hbb06cae1),
	.w3(32'h3ba33d70),
	.w4(32'hbbd87911),
	.w5(32'h3b8a581a),
	.w6(32'hba853d40),
	.w7(32'h3bc8db3b),
	.w8(32'h3ad7173e),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3879151d),
	.w1(32'hbc69de7b),
	.w2(32'h3c1a5ba0),
	.w3(32'hbb937b1a),
	.w4(32'h3c4cf476),
	.w5(32'hbccbe954),
	.w6(32'h3b0207b4),
	.w7(32'h3cd03760),
	.w8(32'hbcb86938),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b03a003),
	.w1(32'h3d19153a),
	.w2(32'hbd683435),
	.w3(32'h3c7706e1),
	.w4(32'h3c5a51b3),
	.w5(32'h3d04ee26),
	.w6(32'hbcb2c0b5),
	.w7(32'hbd0f7243),
	.w8(32'h3d8bf9de),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cfa2289),
	.w1(32'h3a397b85),
	.w2(32'h3ae27a52),
	.w3(32'hbd121527),
	.w4(32'hbb247d22),
	.w5(32'hbacc3a91),
	.w6(32'hbc90af96),
	.w7(32'hbba7ea0c),
	.w8(32'hbae34f64),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8743a1f),
	.w1(32'hbc0d459d),
	.w2(32'hbc311f51),
	.w3(32'h39a16b61),
	.w4(32'hbaff4552),
	.w5(32'hbb1f3f95),
	.w6(32'hbb0f975b),
	.w7(32'h3b30656b),
	.w8(32'hbc3bb947),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb89b70c),
	.w1(32'hbaf127a4),
	.w2(32'h3b81427f),
	.w3(32'hbcf2daf6),
	.w4(32'hbbb4190a),
	.w5(32'hbb828fe5),
	.w6(32'h3c715513),
	.w7(32'h3b14aff7),
	.w8(32'h3c59c6d7),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf15721),
	.w1(32'hbb01f85f),
	.w2(32'h3b5b0719),
	.w3(32'h3be1560d),
	.w4(32'h39def8e9),
	.w5(32'h3b375434),
	.w6(32'hb9f5f1ec),
	.w7(32'hb9ba1370),
	.w8(32'hb85cb716),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b118ca7),
	.w1(32'hbcde7a8c),
	.w2(32'h3b9c93eb),
	.w3(32'hbaa53141),
	.w4(32'hbc2c996b),
	.w5(32'hbc2e8701),
	.w6(32'hba9ada2e),
	.w7(32'hbb50a332),
	.w8(32'hbc48f3df),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc488110),
	.w1(32'hbbf42303),
	.w2(32'h3aada8e6),
	.w3(32'h3b452a0f),
	.w4(32'hba9ae755),
	.w5(32'h3ba395fe),
	.w6(32'hbca5dccd),
	.w7(32'hba950e7e),
	.w8(32'hbaee68cd),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf697fd),
	.w1(32'h3b22d8af),
	.w2(32'h3bbf0d98),
	.w3(32'hbb00f538),
	.w4(32'h391b3cea),
	.w5(32'h3b54d0d3),
	.w6(32'h3b7e3773),
	.w7(32'h3a46a526),
	.w8(32'h3a149c1f),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabec902),
	.w1(32'h3b1ee6ad),
	.w2(32'h3b0b07c5),
	.w3(32'h3af08f94),
	.w4(32'h3c124a13),
	.w5(32'h3b9f617f),
	.w6(32'h3bb46087),
	.w7(32'h3ae28276),
	.w8(32'h3b80da23),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc462148),
	.w1(32'hbb1af873),
	.w2(32'hb9ed199e),
	.w3(32'h3b2c8316),
	.w4(32'hbc0c2b21),
	.w5(32'hba8023f2),
	.w6(32'hbad70aed),
	.w7(32'hbb960d43),
	.w8(32'hbbd9546a),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2a2484),
	.w1(32'hb9bccedd),
	.w2(32'h3b40cd8a),
	.w3(32'hbb68db98),
	.w4(32'hba2158b4),
	.w5(32'h39a0d2b2),
	.w6(32'hbadfd72c),
	.w7(32'hb9c179ea),
	.w8(32'h3a13f1c1),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8432b0),
	.w1(32'h3cc39c0e),
	.w2(32'hbc9eeb54),
	.w3(32'h3a4901b4),
	.w4(32'hbc244107),
	.w5(32'h3bafb23b),
	.w6(32'hbabcc18a),
	.w7(32'hbcbace9f),
	.w8(32'h3c9fc1be),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd79796),
	.w1(32'hba355aeb),
	.w2(32'hbb34e029),
	.w3(32'hbae01c5f),
	.w4(32'h3ac182a9),
	.w5(32'hbad19800),
	.w6(32'hbbd23831),
	.w7(32'h3b5c1fb0),
	.w8(32'hba8ec951),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2ba1dd),
	.w1(32'h3b50c5c5),
	.w2(32'hbbbc3959),
	.w3(32'hbb03add8),
	.w4(32'h3b9b34a9),
	.w5(32'h3b248b27),
	.w6(32'h3b02b47a),
	.w7(32'hbaf97bb4),
	.w8(32'h3aaf7406),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb187142),
	.w1(32'hbca825e3),
	.w2(32'h3c0b4f10),
	.w3(32'h36aacc44),
	.w4(32'h3b234cff),
	.w5(32'hbc6499d6),
	.w6(32'h3b9178b1),
	.w7(32'h3bd55619),
	.w8(32'hbb5bd2e0),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbeb47c),
	.w1(32'h3bf0b883),
	.w2(32'h3c99b000),
	.w3(32'h3cd2229c),
	.w4(32'hbd06b180),
	.w5(32'h3cd23b0a),
	.w6(32'hbbec40ae),
	.w7(32'hbc83a545),
	.w8(32'hbc990b78),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc10fde4),
	.w1(32'hbb23a998),
	.w2(32'h3b094a14),
	.w3(32'hbc3c9362),
	.w4(32'hbb3912e2),
	.w5(32'hbc51f5ce),
	.w6(32'h3ccdca4b),
	.w7(32'hbba5c7e2),
	.w8(32'hbc6293d6),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb185e3c),
	.w1(32'hbbb769b1),
	.w2(32'hbc073059),
	.w3(32'hbc8cd164),
	.w4(32'hbbf2b404),
	.w5(32'hb99fec12),
	.w6(32'hbc1a031c),
	.w7(32'hbbdf95c6),
	.w8(32'h3aa52853),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb649cc4),
	.w1(32'h3b545b18),
	.w2(32'h3b9e3cfe),
	.w3(32'h3c352980),
	.w4(32'hba070151),
	.w5(32'hbae590ab),
	.w6(32'hbc2a1b5f),
	.w7(32'h3c1e48bf),
	.w8(32'h3b218002),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a975f65),
	.w1(32'hbb194af2),
	.w2(32'hbafdec8a),
	.w3(32'h3b924918),
	.w4(32'hbaa9373d),
	.w5(32'h3b02d28b),
	.w6(32'hba8333f3),
	.w7(32'h3af423a8),
	.w8(32'h3b612356),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae2e43b),
	.w1(32'h3b6fc742),
	.w2(32'h3b359e38),
	.w3(32'hbaa1df17),
	.w4(32'h3b1257b8),
	.w5(32'h3b84f0cb),
	.w6(32'h3b051c7e),
	.w7(32'hb99db986),
	.w8(32'h3b3ebbc8),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90d3a2e),
	.w1(32'h3a9134d1),
	.w2(32'h3c07424f),
	.w3(32'h3a4b1387),
	.w4(32'h3bfebc5f),
	.w5(32'h3d044168),
	.w6(32'h3b417209),
	.w7(32'h3c8286f6),
	.w8(32'h3cb1dcaa),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c07e377),
	.w1(32'hbc1dcace),
	.w2(32'hbd131e91),
	.w3(32'h39603107),
	.w4(32'h3c87dcba),
	.w5(32'hbcb92179),
	.w6(32'h3c8477b7),
	.w7(32'hb98abe4b),
	.w8(32'h3cca8b2a),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd047f9),
	.w1(32'hb809755f),
	.w2(32'hbbcdd42a),
	.w3(32'h3adf24cf),
	.w4(32'hb95082c5),
	.w5(32'h3b1690f2),
	.w6(32'hbc4ac97e),
	.w7(32'hbbe22ae8),
	.w8(32'h3c159f8c),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b463458),
	.w1(32'hbb94a40c),
	.w2(32'h3cb1afdf),
	.w3(32'hbbd87b93),
	.w4(32'hbca2bc6e),
	.w5(32'h3c84a828),
	.w6(32'hbbf19cd4),
	.w7(32'h3bdb4e12),
	.w8(32'hbcd960cb),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc647be),
	.w1(32'h3cfeb91c),
	.w2(32'h3d0dd309),
	.w3(32'hbb58077a),
	.w4(32'h3c8710f3),
	.w5(32'h3cb23d08),
	.w6(32'h3cc89ac5),
	.w7(32'h3c7077cb),
	.w8(32'h3d2aafa8),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae5d1ca),
	.w1(32'h3b79d66e),
	.w2(32'h3ba5cbad),
	.w3(32'h3d7d60ee),
	.w4(32'h3bb8416b),
	.w5(32'hb992d426),
	.w6(32'h3c4a1446),
	.w7(32'hbb4685fa),
	.w8(32'hbacf021a),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3d6c8f),
	.w1(32'hbb1d89f8),
	.w2(32'h3bc1fa22),
	.w3(32'h3b96266d),
	.w4(32'hbc168ff6),
	.w5(32'hbb7467a4),
	.w6(32'hba7f0141),
	.w7(32'hb9a7c120),
	.w8(32'hbc04b58c),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb22529f),
	.w1(32'hbbeed9f5),
	.w2(32'h3b771e02),
	.w3(32'h3c37ab3c),
	.w4(32'hbaa9dca4),
	.w5(32'hbbc5e0c0),
	.w6(32'h3c06f4bf),
	.w7(32'hbbe88b09),
	.w8(32'h3ae919ea),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1822d1),
	.w1(32'h3acc5d53),
	.w2(32'hba5199e2),
	.w3(32'h3bbda5bf),
	.w4(32'h3b2d82dc),
	.w5(32'hb83891c6),
	.w6(32'hbb4030e7),
	.w7(32'h3b04285f),
	.w8(32'h3b8ea5f2),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ada0e76),
	.w1(32'h3c2634ae),
	.w2(32'hba2f3d5c),
	.w3(32'hb96d0751),
	.w4(32'hbbfeb3d1),
	.w5(32'hb91b31a8),
	.w6(32'hbb23d5c0),
	.w7(32'hbc7a23fe),
	.w8(32'h3c11652f),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4eeebc),
	.w1(32'h3d43d2bf),
	.w2(32'hbd4d5cf6),
	.w3(32'hbc03f68c),
	.w4(32'hbb58eeee),
	.w5(32'h3d7e89d4),
	.w6(32'hbc3c4775),
	.w7(32'hbd546c6b),
	.w8(32'h3d3300b4),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc5d465),
	.w1(32'hbb65d6fb),
	.w2(32'hbc8eb041),
	.w3(32'hbd9f720e),
	.w4(32'h3cc59480),
	.w5(32'hbd118438),
	.w6(32'h3c6bcfc8),
	.w7(32'h3a6264de),
	.w8(32'h3cc7ac13),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1324ff),
	.w1(32'hba284100),
	.w2(32'h3b05b51d),
	.w3(32'h3c14930a),
	.w4(32'h3a08d2ee),
	.w5(32'h3aed501b),
	.w6(32'hbd25df19),
	.w7(32'h3b54f66e),
	.w8(32'hb879ae02),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba323539),
	.w1(32'h3aaa53a9),
	.w2(32'h3b8e290b),
	.w3(32'hb9667aaf),
	.w4(32'h3b1e2fbb),
	.w5(32'hbb40dd1b),
	.w6(32'h3aee7ccd),
	.w7(32'hbbd00276),
	.w8(32'h3a5c56a4),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8b34ab),
	.w1(32'h3ae9421d),
	.w2(32'hbaca2ce5),
	.w3(32'h3b27190f),
	.w4(32'hbb3942d1),
	.w5(32'hbb6c35e4),
	.w6(32'hbbe2ef87),
	.w7(32'h3b55687f),
	.w8(32'h3ae777ea),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb579891),
	.w1(32'hb9e8dfd1),
	.w2(32'hbaaebd3b),
	.w3(32'hbbed9306),
	.w4(32'hbb021788),
	.w5(32'hbbb7970d),
	.w6(32'hbb0782e8),
	.w7(32'hbaa48b40),
	.w8(32'hbb5322ad),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4cf348),
	.w1(32'hbc93da4d),
	.w2(32'hbb127116),
	.w3(32'hbb142456),
	.w4(32'h3b1fcac9),
	.w5(32'hbccaa88c),
	.w6(32'hbb54c2e5),
	.w7(32'h3cbef892),
	.w8(32'hbcdb5ded),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7cb7c8),
	.w1(32'hbc23d950),
	.w2(32'hbc061881),
	.w3(32'hbc4309a3),
	.w4(32'h3ac5ffac),
	.w5(32'hbadb5dce),
	.w6(32'h3c03b5d1),
	.w7(32'h3b09400b),
	.w8(32'hbc2cefb8),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb079efc),
	.w1(32'hbbe53924),
	.w2(32'hbca9e4d3),
	.w3(32'hbbbf9a99),
	.w4(32'hbc500d1c),
	.w5(32'hbbf7f7b9),
	.w6(32'h3bc813c3),
	.w7(32'hbcb20dfb),
	.w8(32'hbc2ca606),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfd858a),
	.w1(32'h39c1d970),
	.w2(32'h3b55a57b),
	.w3(32'hbaba53cd),
	.w4(32'hba5dfc98),
	.w5(32'hb5a58aea),
	.w6(32'h3b395fa7),
	.w7(32'h3adb60b1),
	.w8(32'hbb1536dd),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bedd4b2),
	.w1(32'hbd1a21c4),
	.w2(32'h3d74fbcb),
	.w3(32'h3b35f578),
	.w4(32'hbc1edda6),
	.w5(32'hbd02df0f),
	.w6(32'hb92f34a5),
	.w7(32'h3d491554),
	.w8(32'hbd94b89e),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule