module layer_8_featuremap_15(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5fa42b),
	.w1(32'h3cd96720),
	.w2(32'h3bf656b2),
	.w3(32'hbc09860b),
	.w4(32'h3d103bf3),
	.w5(32'hbc9e1bbe),
	.w6(32'hbb7c7eff),
	.w7(32'hbca3e2f0),
	.w8(32'h3c9b304c),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc961122),
	.w1(32'h3ae47d02),
	.w2(32'hbc023606),
	.w3(32'hbb631008),
	.w4(32'hbbb8e446),
	.w5(32'hbc3440aa),
	.w6(32'hbcd52d59),
	.w7(32'hbd223145),
	.w8(32'h3bd1e1f8),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4c0511),
	.w1(32'hbc3e3196),
	.w2(32'hbc8b8c27),
	.w3(32'hbc5fd373),
	.w4(32'hbad3400d),
	.w5(32'hbcdeda3c),
	.w6(32'hbadb5496),
	.w7(32'h39b7fd32),
	.w8(32'h3bea082e),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d497e29),
	.w1(32'hbceec8e8),
	.w2(32'hbb19d6df),
	.w3(32'h3b3fe4bc),
	.w4(32'hbbe088ec),
	.w5(32'h3af24383),
	.w6(32'h3c100b50),
	.w7(32'hbcac9c8e),
	.w8(32'hbb4724c8),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb2a410),
	.w1(32'h3c93788c),
	.w2(32'hbc8d708d),
	.w3(32'hb9811f94),
	.w4(32'hb94acb3d),
	.w5(32'hba9a82ae),
	.w6(32'hbc85aa20),
	.w7(32'h3c4bdc9d),
	.w8(32'h3a975e29),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe56652),
	.w1(32'hbbf07452),
	.w2(32'hbc69e367),
	.w3(32'hbca841b5),
	.w4(32'hbbd07522),
	.w5(32'hbca40522),
	.w6(32'hbb7bc309),
	.w7(32'hbb0fbabf),
	.w8(32'hb950458e),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc90657f),
	.w1(32'hbc215f9a),
	.w2(32'h3a44ed49),
	.w3(32'hbc472e38),
	.w4(32'hbbfb01da),
	.w5(32'hbc5a53db),
	.w6(32'h3d0bc68f),
	.w7(32'hbb8bf4eb),
	.w8(32'hbb097e38),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd411e9),
	.w1(32'hbc155de4),
	.w2(32'h3cac7b27),
	.w3(32'h3a74e15f),
	.w4(32'h3c703a15),
	.w5(32'hbbb17ee1),
	.w6(32'h3d043991),
	.w7(32'h3d68c9fa),
	.w8(32'hbb2656c2),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b96fc68),
	.w1(32'hbc60610c),
	.w2(32'hbc42b069),
	.w3(32'hbb7103c5),
	.w4(32'hbb51e9c0),
	.w5(32'hbb82c0ca),
	.w6(32'h3b4f7071),
	.w7(32'hbab6f99d),
	.w8(32'hbbbb580d),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbfcd7d),
	.w1(32'hbc361ded),
	.w2(32'hbc70c15d),
	.w3(32'h3d3bad55),
	.w4(32'h3d0ee8a2),
	.w5(32'hbc18999c),
	.w6(32'hbc454db3),
	.w7(32'h3d4ab943),
	.w8(32'h3b74a4d2),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d0f303e),
	.w1(32'h3abe3b9b),
	.w2(32'h3c471b66),
	.w3(32'hbc9e99be),
	.w4(32'hbc7cbf65),
	.w5(32'hbc48d7cd),
	.w6(32'hbc07172c),
	.w7(32'hbc1cbbd9),
	.w8(32'h3b74861a),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb0d488),
	.w1(32'hbcaa0307),
	.w2(32'h3c2629ab),
	.w3(32'h3c10c0db),
	.w4(32'h3acd8735),
	.w5(32'h39aa0de6),
	.w6(32'hbb83b73d),
	.w7(32'hbc96128d),
	.w8(32'h3d3d438d),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb08085a),
	.w1(32'hbc2721cd),
	.w2(32'hbc112f60),
	.w3(32'h3c0527da),
	.w4(32'h3b4f65b2),
	.w5(32'hba3b4135),
	.w6(32'hbbd75185),
	.w7(32'hbc3ee318),
	.w8(32'hbb93b8bf),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb83f702),
	.w1(32'hbc903b60),
	.w2(32'hbc40ba0c),
	.w3(32'hbcbfd04b),
	.w4(32'hba4c2223),
	.w5(32'h3bcdc025),
	.w6(32'hbbd611be),
	.w7(32'hbd27ed61),
	.w8(32'h3bf2c644),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc721395),
	.w1(32'h3b568489),
	.w2(32'hbcbe2c50),
	.w3(32'hbb4878e1),
	.w4(32'h3af8d015),
	.w5(32'hbc37b787),
	.w6(32'hbb910914),
	.w7(32'h3a394602),
	.w8(32'h3a96c0f1),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b214ab5),
	.w1(32'h3c2bf505),
	.w2(32'h3c006fc1),
	.w3(32'hbc030b0d),
	.w4(32'hbbfa9281),
	.w5(32'h3d047b37),
	.w6(32'h3b14b55f),
	.w7(32'hba548001),
	.w8(32'h3a4d0879),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8b25fa),
	.w1(32'hbb042e22),
	.w2(32'h388366f2),
	.w3(32'h3c5a2cc3),
	.w4(32'hba478fd2),
	.w5(32'hbc00cf6d),
	.w6(32'h3a45508d),
	.w7(32'hbbd0b80d),
	.w8(32'h3b927415),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e3dbbb),
	.w1(32'h3b12c71f),
	.w2(32'hbc1fc72c),
	.w3(32'h3cedf33b),
	.w4(32'h398e4966),
	.w5(32'hbc703fc8),
	.w6(32'h3ce6f8ba),
	.w7(32'hbc56e4d0),
	.w8(32'h39f00b22),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd4b0d80),
	.w1(32'h3baec363),
	.w2(32'h3cfcca76),
	.w3(32'hbc53cbf8),
	.w4(32'hba7f24e8),
	.w5(32'h3cd4e91c),
	.w6(32'h3b3e6cae),
	.w7(32'hbcc0185e),
	.w8(32'hbcb726d6),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac1d5b0),
	.w1(32'hbce25f56),
	.w2(32'h3ce2607e),
	.w3(32'h3c2ec314),
	.w4(32'hbcc0b6df),
	.w5(32'h3c4b93bc),
	.w6(32'hbb3533df),
	.w7(32'h3d072e18),
	.w8(32'h3b9beb75),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c157121),
	.w1(32'hbbd31a6c),
	.w2(32'h3b5b16f3),
	.w3(32'hb9e23b72),
	.w4(32'hbcae1a6c),
	.w5(32'hbb017a40),
	.w6(32'h3c423afc),
	.w7(32'h3ad7b7fe),
	.w8(32'hbb445bbb),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa57103),
	.w1(32'hbb22fdaa),
	.w2(32'hbbc02dab),
	.w3(32'h3bef6aed),
	.w4(32'h3adc0363),
	.w5(32'hbbc51ccf),
	.w6(32'h3c439edf),
	.w7(32'h3c34be5d),
	.w8(32'h3986a10c),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0effc1),
	.w1(32'h3cd49903),
	.w2(32'h3c3ce2dd),
	.w3(32'hbca23c1c),
	.w4(32'hbbb0448d),
	.w5(32'h3c3d7997),
	.w6(32'hbc7eda71),
	.w7(32'hbc3574b8),
	.w8(32'h3b5961a2),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b69f3d5),
	.w1(32'hbc04f286),
	.w2(32'hbc19b831),
	.w3(32'hbc8b6600),
	.w4(32'hb6885fe8),
	.w5(32'h3abe2f13),
	.w6(32'hba3e23ed),
	.w7(32'h3aa6e9a9),
	.w8(32'h3b4834b1),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf008ec),
	.w1(32'h3c8c110b),
	.w2(32'h3b4ac6ff),
	.w3(32'h3b85afc9),
	.w4(32'h3b214c35),
	.w5(32'h3be14288),
	.w6(32'h3aa9f0dc),
	.w7(32'hb9ff3273),
	.w8(32'hbb22818c),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba38b7a1),
	.w1(32'h3c22acce),
	.w2(32'h3be9b14c),
	.w3(32'hbc78cd5d),
	.w4(32'h3bff6bf3),
	.w5(32'h3aeb6dd7),
	.w6(32'hbc76720f),
	.w7(32'hbabcb8e1),
	.w8(32'h3abca224),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad811ab),
	.w1(32'hbc020be0),
	.w2(32'hbb6b8ade),
	.w3(32'hbbc98b24),
	.w4(32'hbbfb95fc),
	.w5(32'h3cd23e20),
	.w6(32'h3bf1a970),
	.w7(32'h3b49ea44),
	.w8(32'hbba97e9e),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd5ec2f8),
	.w1(32'hbd19ea63),
	.w2(32'h3df0f9e5),
	.w3(32'hbd3456af),
	.w4(32'hbd812f6c),
	.w5(32'hbbdc03cc),
	.w6(32'h3d28f888),
	.w7(32'hbd1a14fc),
	.w8(32'hbd767b78),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3f4298),
	.w1(32'hbb47f64a),
	.w2(32'h3c9d0933),
	.w3(32'h3b70fde7),
	.w4(32'h3c2ddb6f),
	.w5(32'hbc5ad846),
	.w6(32'hbcbbb163),
	.w7(32'h3c003faf),
	.w8(32'hbd3ff97e),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf97b71),
	.w1(32'hbce5e432),
	.w2(32'hbd399bef),
	.w3(32'hbcf099ba),
	.w4(32'h3b9b4850),
	.w5(32'hba52209a),
	.w6(32'hbc166bc1),
	.w7(32'hbbca0960),
	.w8(32'h3c93a3af),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca1a505),
	.w1(32'hbca9f577),
	.w2(32'hbbb3595b),
	.w3(32'hbbab54a3),
	.w4(32'hbc1e9d62),
	.w5(32'hbbf5c8bc),
	.w6(32'hbac6acd1),
	.w7(32'hbc1d058c),
	.w8(32'h3b435d33),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9133ac),
	.w1(32'hbb8f614b),
	.w2(32'h3ad8ebbe),
	.w3(32'h3b6fb3cc),
	.w4(32'hbd0f4c0f),
	.w5(32'hbc9d9e05),
	.w6(32'hbbfccad1),
	.w7(32'h3c98cd7e),
	.w8(32'hbc8b25fa),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fa0a35),
	.w1(32'hbb43c85c),
	.w2(32'hbc26a69f),
	.w3(32'hbc502dd0),
	.w4(32'hbc72aa06),
	.w5(32'h3d0938e9),
	.w6(32'hbc725aac),
	.w7(32'hba173b44),
	.w8(32'hbcaef8b7),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb7c35a),
	.w1(32'hbb57dab9),
	.w2(32'hbb251a7f),
	.w3(32'h3d92d045),
	.w4(32'hbc7001fe),
	.w5(32'h3c18d1db),
	.w6(32'h3addff35),
	.w7(32'hbcff0c3a),
	.w8(32'hbbbb0ff5),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c39a6ac),
	.w1(32'hbd0dc5ec),
	.w2(32'hbd174eb4),
	.w3(32'hbbfce53b),
	.w4(32'hbd0721ce),
	.w5(32'hbc8f1386),
	.w6(32'hb9b30ab0),
	.w7(32'hbcb0b877),
	.w8(32'hbc0152dd),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4f896a),
	.w1(32'hbc049e0c),
	.w2(32'h3c0f740a),
	.w3(32'hbbad55fa),
	.w4(32'h3cb4cb22),
	.w5(32'hbcc9c285),
	.w6(32'h3d57af92),
	.w7(32'hbb984828),
	.w8(32'hbc9e8196),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b50b651),
	.w1(32'hbc4678ba),
	.w2(32'h395db8c2),
	.w3(32'h3ba67680),
	.w4(32'hb9ac561e),
	.w5(32'hbc5823b5),
	.w6(32'hbce1f940),
	.w7(32'h3b760320),
	.w8(32'hbb4dabc3),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc37a9ed),
	.w1(32'h3cb36054),
	.w2(32'h3c796fdd),
	.w3(32'h3a089333),
	.w4(32'h3a6685f2),
	.w5(32'h3c980078),
	.w6(32'h3b977ae0),
	.w7(32'h3bfb5839),
	.w8(32'h3c77bca0),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc877842),
	.w1(32'hbbb81ddc),
	.w2(32'h3b7a857a),
	.w3(32'hbcb187c7),
	.w4(32'h3cde76d1),
	.w5(32'h3b328dd9),
	.w6(32'hbc267733),
	.w7(32'hbbafec39),
	.w8(32'h3c845802),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc076aa),
	.w1(32'h3c809e10),
	.w2(32'hbbc03d39),
	.w3(32'h3b3de969),
	.w4(32'hba3c2a86),
	.w5(32'hbc49ef98),
	.w6(32'hbc3098a8),
	.w7(32'hbc292823),
	.w8(32'h3c82c4e0),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdb77b9),
	.w1(32'h3c9f6a9b),
	.w2(32'h3cd75396),
	.w3(32'h3c0d5f8a),
	.w4(32'h3c23e478),
	.w5(32'h3c55de90),
	.w6(32'hbd079d49),
	.w7(32'hbae902b3),
	.w8(32'h3c537cc8),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a2f151),
	.w1(32'hbc105f4d),
	.w2(32'h3c2c5c65),
	.w3(32'hbb5ff5c3),
	.w4(32'h3c6d1b50),
	.w5(32'hbc46d929),
	.w6(32'hbb1b2f01),
	.w7(32'hbbc09b52),
	.w8(32'hbbcde740),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1ea62f),
	.w1(32'hbb168ecf),
	.w2(32'hbc1159d5),
	.w3(32'hbc5ed722),
	.w4(32'hbc91d6ae),
	.w5(32'hbbe5f9db),
	.w6(32'hbb850cd7),
	.w7(32'hbad2de52),
	.w8(32'hbc97567e),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4fe444),
	.w1(32'h3d77be34),
	.w2(32'h3c3ffe3c),
	.w3(32'hbca7c628),
	.w4(32'hbcb9dbc4),
	.w5(32'hbb266727),
	.w6(32'hbb233c9b),
	.w7(32'hbbadb26a),
	.w8(32'h3d342a4b),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8cef9e),
	.w1(32'h3cff0f7a),
	.w2(32'hba0ee5c5),
	.w3(32'h3c89aa2b),
	.w4(32'h3ae884ff),
	.w5(32'h3cd40400),
	.w6(32'hbc377399),
	.w7(32'hbc093b8c),
	.w8(32'h3c61cd65),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc687a1e),
	.w1(32'hbb413ddf),
	.w2(32'h3b1f9a77),
	.w3(32'hbb5ce282),
	.w4(32'hbb27bdf2),
	.w5(32'h3c013798),
	.w6(32'h3b6a9e40),
	.w7(32'hbb909c29),
	.w8(32'hbbbce1f9),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9fd4cc),
	.w1(32'hbc4d82fb),
	.w2(32'hbbe3d622),
	.w3(32'hbbb81692),
	.w4(32'hbc586ad5),
	.w5(32'hbc6daf19),
	.w6(32'hbd0ef207),
	.w7(32'h3d252d86),
	.w8(32'hbbad3e32),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37abb162),
	.w1(32'hbcc5cdce),
	.w2(32'h3ba069a8),
	.w3(32'h3c5b9807),
	.w4(32'h3b021c94),
	.w5(32'h3be4079b),
	.w6(32'hbb1b989c),
	.w7(32'h39a04514),
	.w8(32'hbc301cdf),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c16a7f6),
	.w1(32'hbba5b5af),
	.w2(32'h3b37ecb6),
	.w3(32'hbc0c1534),
	.w4(32'hbc81c690),
	.w5(32'hbc758970),
	.w6(32'hbb3650d3),
	.w7(32'h3da65db4),
	.w8(32'hbb136a2f),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0b07dd),
	.w1(32'h3bcebcee),
	.w2(32'h3b6a2ed3),
	.w3(32'hbc749c4b),
	.w4(32'h3b2b8b81),
	.w5(32'h3bec8469),
	.w6(32'h3d3b8389),
	.w7(32'hbbce8196),
	.w8(32'h3b56bc9a),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d10120e),
	.w1(32'h3d0678e9),
	.w2(32'h3be13deb),
	.w3(32'h3bd21538),
	.w4(32'h3c07bbe0),
	.w5(32'h3c3391fb),
	.w6(32'h3c3b7ad2),
	.w7(32'h3c25fb57),
	.w8(32'h3a7dc879),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcdb1111),
	.w1(32'h3ccd4d53),
	.w2(32'h3cd6bd8b),
	.w3(32'hbc443ea6),
	.w4(32'h3a7a7e52),
	.w5(32'h3d999e8d),
	.w6(32'hbc96559c),
	.w7(32'hbc0cc734),
	.w8(32'h3ccc8791),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6cdc2d),
	.w1(32'hbb12f46f),
	.w2(32'h3cfe560b),
	.w3(32'hbd0e10b8),
	.w4(32'h3aba9d08),
	.w5(32'h3ca88990),
	.w6(32'h3d07c186),
	.w7(32'h3c2506bd),
	.w8(32'hbb07020f),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0e2044),
	.w1(32'hbc15c900),
	.w2(32'h3bcd5de8),
	.w3(32'h3d0f2e55),
	.w4(32'h3c08513d),
	.w5(32'hba9d5f42),
	.w6(32'hbae5c5c1),
	.w7(32'hbbe96bf9),
	.w8(32'hba1272fc),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb829b73),
	.w1(32'h3acb199f),
	.w2(32'hb9848624),
	.w3(32'hbb987887),
	.w4(32'hbc3b18c1),
	.w5(32'hbc2230bf),
	.w6(32'h3c00e1a9),
	.w7(32'h3a15e5a2),
	.w8(32'hbc1964cb),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0d5263),
	.w1(32'hbbf43c7b),
	.w2(32'h3d328316),
	.w3(32'h3cbd409f),
	.w4(32'h3c3d55db),
	.w5(32'h3c69ee27),
	.w6(32'hbc8d0fa2),
	.w7(32'hbc41f94f),
	.w8(32'h3d115438),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc79add),
	.w1(32'hbc3973a5),
	.w2(32'hbc299c7f),
	.w3(32'h3b65e3cc),
	.w4(32'hbb9e3e53),
	.w5(32'hbb64541d),
	.w6(32'h3b8a166b),
	.w7(32'h3b0e7194),
	.w8(32'h3b3a37b9),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c96590a),
	.w1(32'h3b653cb7),
	.w2(32'h3ca980b9),
	.w3(32'hbb13ddb9),
	.w4(32'h3abee169),
	.w5(32'h3cc49354),
	.w6(32'h3b484207),
	.w7(32'hbc4d4e4e),
	.w8(32'h3b974ffc),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb72d55a),
	.w1(32'hbc0b4c71),
	.w2(32'h3bf832f3),
	.w3(32'hbc40fa7b),
	.w4(32'hbb76ca8e),
	.w5(32'hbbb5fbd7),
	.w6(32'h3c97f9a3),
	.w7(32'h3c4c27f5),
	.w8(32'h390bd8f8),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c49da5e),
	.w1(32'h3c50275b),
	.w2(32'h3caccfab),
	.w3(32'h3c3cde69),
	.w4(32'h3c3f68f6),
	.w5(32'h3c01b79e),
	.w6(32'h3b84fdb1),
	.w7(32'h3c15054b),
	.w8(32'h3c803bd5),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a52fdbf),
	.w1(32'h3b660f38),
	.w2(32'h3cc24271),
	.w3(32'h3bba3813),
	.w4(32'hbcdee05d),
	.w5(32'hbb0234cd),
	.w6(32'hba876493),
	.w7(32'h3a4d3d43),
	.w8(32'hbbc079f4),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc77cf7),
	.w1(32'h3cbff074),
	.w2(32'h3b2341e8),
	.w3(32'hbc0b1ceb),
	.w4(32'hbc687705),
	.w5(32'hba639954),
	.w6(32'hbc0d1dd4),
	.w7(32'hbb0d60be),
	.w8(32'h3cc543ed),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb11baa0),
	.w1(32'h3ba63955),
	.w2(32'h3d85b182),
	.w3(32'h3c36db7d),
	.w4(32'h3c2726a1),
	.w5(32'h3b1642dd),
	.w6(32'hbc1c70a7),
	.w7(32'h3c166a4c),
	.w8(32'hbb5b321f),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c081676),
	.w1(32'h3bccdc07),
	.w2(32'h3c36ef2f),
	.w3(32'h3b46a865),
	.w4(32'h3d024f18),
	.w5(32'h3a105d11),
	.w6(32'hbbe645a9),
	.w7(32'h3b571339),
	.w8(32'h3a89e33a),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0284e6),
	.w1(32'hbbd4c9ee),
	.w2(32'hbb987119),
	.w3(32'hbc2c1d17),
	.w4(32'h3b350017),
	.w5(32'hbb016656),
	.w6(32'hba115713),
	.w7(32'h3d5e4323),
	.w8(32'hba5ac7b7),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb30c742),
	.w1(32'hbb04dcd6),
	.w2(32'hbb59f24d),
	.w3(32'hbb824f29),
	.w4(32'hbbdc65dd),
	.w5(32'h3bb76155),
	.w6(32'h3b37d89d),
	.w7(32'hba879562),
	.w8(32'hbb328ed6),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a209473),
	.w1(32'hbb23f372),
	.w2(32'hbb8d6455),
	.w3(32'h3c7bcccc),
	.w4(32'hbc563d54),
	.w5(32'hbbce097e),
	.w6(32'h3bb45a2e),
	.w7(32'h3b9ef8ff),
	.w8(32'h3b0370d3),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc11666e),
	.w1(32'h3b120948),
	.w2(32'h3b82bbce),
	.w3(32'h3c0c933d),
	.w4(32'hbb890a33),
	.w5(32'h3b2cb124),
	.w6(32'hbb85e84f),
	.w7(32'hbc5058cb),
	.w8(32'hbb989ce6),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3148f2),
	.w1(32'hbb0c291b),
	.w2(32'hbc42e4bd),
	.w3(32'hbb96b43d),
	.w4(32'h3c6aaef8),
	.w5(32'h3b5036d9),
	.w6(32'hbc34dc07),
	.w7(32'hb97dd58a),
	.w8(32'hbb01d7a3),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc37a850),
	.w1(32'hbbbab2cf),
	.w2(32'h3cb89997),
	.w3(32'hbc330cf9),
	.w4(32'hbb281644),
	.w5(32'h3b330c9a),
	.w6(32'h3bf56811),
	.w7(32'hbbeb1fba),
	.w8(32'h3d2cac9c),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfd9367),
	.w1(32'h3c521787),
	.w2(32'hbc9891cc),
	.w3(32'h3cd472d1),
	.w4(32'h398c3599),
	.w5(32'h3cb8cd52),
	.w6(32'hbc051a4b),
	.w7(32'hbce0d4b8),
	.w8(32'hbc976281),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb351a21),
	.w1(32'h3a999518),
	.w2(32'h3bc79120),
	.w3(32'h3be00df6),
	.w4(32'h3c436aed),
	.w5(32'hbc8a45f0),
	.w6(32'hbbae667e),
	.w7(32'hbc918d77),
	.w8(32'hbd0bc0e0),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2fc215),
	.w1(32'hbc83e69f),
	.w2(32'h3c4fe5b2),
	.w3(32'hbd03e223),
	.w4(32'hb9847835),
	.w5(32'hbc2466f7),
	.w6(32'h3af78470),
	.w7(32'h3d711356),
	.w8(32'h3a868228),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4fd719),
	.w1(32'hbbfd13c5),
	.w2(32'h3cd48b0d),
	.w3(32'h3c8afa43),
	.w4(32'hbc8fad21),
	.w5(32'hbd07d954),
	.w6(32'h3c9fe08e),
	.w7(32'h3bee03f4),
	.w8(32'hbbcaebf9),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab22ef4),
	.w1(32'h3c69a704),
	.w2(32'hbc2b4b3b),
	.w3(32'hbc93a217),
	.w4(32'hbc564e34),
	.w5(32'hbc19dc77),
	.w6(32'h3c76d6c1),
	.w7(32'hbbb045f9),
	.w8(32'hbbb85c81),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d0e7d91),
	.w1(32'hbb8cdf07),
	.w2(32'h3cd8d47c),
	.w3(32'hbc0318d9),
	.w4(32'h3c6b4d1a),
	.w5(32'h3d412da9),
	.w6(32'hbc13388f),
	.w7(32'h3b21ee49),
	.w8(32'h3ae6892b),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9ee31f),
	.w1(32'h3b6fed0c),
	.w2(32'h3bae74f0),
	.w3(32'hbc979ad4),
	.w4(32'hbbc6bf4c),
	.w5(32'hbc7d2eea),
	.w6(32'h3b367e1d),
	.w7(32'h3c3c6744),
	.w8(32'h3c9aa1d7),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd56f81),
	.w1(32'hbc731ce1),
	.w2(32'h3bff6a1e),
	.w3(32'h3c8c6cc3),
	.w4(32'h3bd2b4bf),
	.w5(32'h3c0390e8),
	.w6(32'hbc67fc74),
	.w7(32'hbbf382d8),
	.w8(32'h3c43d775),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb96d67c),
	.w1(32'h3c9e137f),
	.w2(32'h3a9e5961),
	.w3(32'h3c5200f2),
	.w4(32'h3b7256b1),
	.w5(32'h3c78b1bc),
	.w6(32'h3af7c9c6),
	.w7(32'hbad26404),
	.w8(32'h3c718834),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7a4637),
	.w1(32'hba30ddaa),
	.w2(32'h3b3cc476),
	.w3(32'hba0f0de8),
	.w4(32'h3a74ed72),
	.w5(32'h3c230776),
	.w6(32'h3c528884),
	.w7(32'hbc522862),
	.w8(32'h3b95487a),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb7d090),
	.w1(32'hbbf1a4cc),
	.w2(32'h3bd897c6),
	.w3(32'h393969a7),
	.w4(32'hbaea2c4b),
	.w5(32'hbc77f788),
	.w6(32'hbcc54291),
	.w7(32'h3c6bb2d1),
	.w8(32'h3bf54de6),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a49ba0b),
	.w1(32'h3c507ef9),
	.w2(32'hbc0baa86),
	.w3(32'h3cdca7ab),
	.w4(32'h3c946e3f),
	.w5(32'h3cc1b3cc),
	.w6(32'hbb1e5e23),
	.w7(32'h3c0d7a93),
	.w8(32'h3c05d37a),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a25424),
	.w1(32'hbc1a2a9d),
	.w2(32'h3d9750b6),
	.w3(32'h3b49283b),
	.w4(32'hbcb8fb3a),
	.w5(32'h3babac16),
	.w6(32'hbc7fc1ce),
	.w7(32'hbb57eb99),
	.w8(32'h3c26ed04),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d8ae6c3),
	.w1(32'h3d4ce127),
	.w2(32'h3d5d5ed6),
	.w3(32'h3d2c9bd9),
	.w4(32'h3c8ea823),
	.w5(32'h3d517c47),
	.w6(32'h3ad557e7),
	.w7(32'hbb862c02),
	.w8(32'h3cc24090),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc809a7b),
	.w1(32'h3c768def),
	.w2(32'h3cf461c9),
	.w3(32'hbc200f5d),
	.w4(32'hbb45d325),
	.w5(32'h3bf3c25a),
	.w6(32'hbc22a333),
	.w7(32'hbc79491a),
	.w8(32'hbc680d9c),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c802d00),
	.w1(32'h3cab8fa5),
	.w2(32'h3cc2f70d),
	.w3(32'h3bbc0253),
	.w4(32'h3c898331),
	.w5(32'h3cd4ec45),
	.w6(32'hbc010261),
	.w7(32'h3b998554),
	.w8(32'h3ca0eff4),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bccd5fd),
	.w1(32'h3b53e30e),
	.w2(32'h3bd2cab6),
	.w3(32'hbae41dd0),
	.w4(32'hb95643f2),
	.w5(32'h3b0174f7),
	.w6(32'h3be12797),
	.w7(32'h3a887d33),
	.w8(32'hbb8744ad),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b74d11b),
	.w1(32'h3a95975b),
	.w2(32'h3a7f96d7),
	.w3(32'hbbc64573),
	.w4(32'h3c01da52),
	.w5(32'h39e9c91f),
	.w6(32'h3beb2ac4),
	.w7(32'h3c18d1a0),
	.w8(32'h3944633d),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb919c815),
	.w1(32'hbbd73aa2),
	.w2(32'h3aebf385),
	.w3(32'h3c1d93ff),
	.w4(32'hba369240),
	.w5(32'h3b0aa505),
	.w6(32'h3a91f781),
	.w7(32'h3936de64),
	.w8(32'hbc6d027c),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb807749),
	.w1(32'h3acda848),
	.w2(32'h3bf29675),
	.w3(32'hbbea749b),
	.w4(32'hbac2062b),
	.w5(32'h3bac6bfc),
	.w6(32'hbb624a47),
	.w7(32'hba9b9cc7),
	.w8(32'hbb5b50dd),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c37690e),
	.w1(32'h3ba18cbc),
	.w2(32'h3ceac81f),
	.w3(32'h3bcc2999),
	.w4(32'h3c63979a),
	.w5(32'h3b8583e1),
	.w6(32'h3b8776d3),
	.w7(32'h3c785254),
	.w8(32'hbb4bf4a5),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8cc959),
	.w1(32'hbaf22f44),
	.w2(32'hbb95ed11),
	.w3(32'h3b8d0d37),
	.w4(32'hbbf1ccad),
	.w5(32'hba4d6a22),
	.w6(32'hbbce0290),
	.w7(32'h3bc9aa96),
	.w8(32'h3bc4df32),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcb18cb),
	.w1(32'hb9e44570),
	.w2(32'hbc1b3279),
	.w3(32'h3b9a5671),
	.w4(32'hb9d34c64),
	.w5(32'hbc22b838),
	.w6(32'h3a9837f6),
	.w7(32'hbb92a76e),
	.w8(32'h3b2c240d),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ecaca4),
	.w1(32'h3a99d24b),
	.w2(32'h3bb21270),
	.w3(32'hbbcb0fa2),
	.w4(32'hbba259a1),
	.w5(32'hbad5852d),
	.w6(32'hba05a921),
	.w7(32'hbb06465b),
	.w8(32'h3c00eb3c),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a3b68),
	.w1(32'hbb033408),
	.w2(32'h3b1130ea),
	.w3(32'hbb9b8bc5),
	.w4(32'h3bb5b5d4),
	.w5(32'h3ba39a0c),
	.w6(32'hbacb8697),
	.w7(32'hbb8bdabb),
	.w8(32'hba8597af),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3dbb1a),
	.w1(32'h3b7046a4),
	.w2(32'h3b6df6bc),
	.w3(32'hbbbce9f3),
	.w4(32'hbb356873),
	.w5(32'h3c22595f),
	.w6(32'hbc1389f7),
	.w7(32'hbbdb953e),
	.w8(32'hbb87f504),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbdb434),
	.w1(32'h3be5ce17),
	.w2(32'h3c830c12),
	.w3(32'hbbff9222),
	.w4(32'h368951ec),
	.w5(32'h3c1cb8c4),
	.w6(32'h3bda230b),
	.w7(32'hbc4228b3),
	.w8(32'hba67a4a2),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1a40bb),
	.w1(32'hbb34d461),
	.w2(32'hbba6371a),
	.w3(32'hbb245464),
	.w4(32'h3c27cf5a),
	.w5(32'hbc33a204),
	.w6(32'hbac196f3),
	.w7(32'hbb6d1ec1),
	.w8(32'h3b3a4b6a),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa5d0fb),
	.w1(32'hbbbf2ba1),
	.w2(32'h3bc9ac1d),
	.w3(32'hbb36351e),
	.w4(32'h3b6d77c4),
	.w5(32'h3b9943aa),
	.w6(32'h3b1aa3fb),
	.w7(32'hbc2ea671),
	.w8(32'hbba4b14c),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c72872d),
	.w1(32'h3b35a421),
	.w2(32'hbaafc75e),
	.w3(32'h3c9f04a9),
	.w4(32'hbb2d955d),
	.w5(32'h3ae73aeb),
	.w6(32'h3add8c44),
	.w7(32'h3b2e9506),
	.w8(32'h3ab95d6f),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c38d966),
	.w1(32'h3c28f5f2),
	.w2(32'h3c61e38c),
	.w3(32'h39c55aea),
	.w4(32'h3c2284f0),
	.w5(32'h3b07a3e4),
	.w6(32'h3ba55770),
	.w7(32'h3b652547),
	.w8(32'hbbc2f0c6),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c37243),
	.w1(32'h3c70e8e4),
	.w2(32'hbb21d509),
	.w3(32'h3aeefcf9),
	.w4(32'h3cad8bf0),
	.w5(32'h3b890cb6),
	.w6(32'hbb874b05),
	.w7(32'h3bb7dae9),
	.w8(32'h3b3d646f),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2e83cb),
	.w1(32'h3ad5ad30),
	.w2(32'h3c229d36),
	.w3(32'hbb3a09d1),
	.w4(32'hbb483210),
	.w5(32'h3b38ca27),
	.w6(32'h3b383362),
	.w7(32'h3b6af067),
	.w8(32'hbc9ed98b),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe74ef0),
	.w1(32'h3c0ba4ff),
	.w2(32'h3c169d70),
	.w3(32'h3cf7371b),
	.w4(32'hbbd17e70),
	.w5(32'hbd803ba3),
	.w6(32'h3c14ed89),
	.w7(32'hbb85f539),
	.w8(32'h3b20ba64),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc82b93),
	.w1(32'hbb123cff),
	.w2(32'h3aafdf97),
	.w3(32'h3be3c4d0),
	.w4(32'hbc85f5df),
	.w5(32'hbb11c185),
	.w6(32'hba910bd7),
	.w7(32'h3bd70073),
	.w8(32'hbc1b6795),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c659dff),
	.w1(32'hbba06203),
	.w2(32'h3cb4c83d),
	.w3(32'h3ad98acd),
	.w4(32'hbc20a461),
	.w5(32'hbaf8eba2),
	.w6(32'hbb4db4d0),
	.w7(32'hbad849cb),
	.w8(32'hbc2d5235),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1bd0c9),
	.w1(32'hbbd487f4),
	.w2(32'h3c4891c6),
	.w3(32'hba9bd9ac),
	.w4(32'h3cf965e3),
	.w5(32'h3c0e1917),
	.w6(32'hbb20dee3),
	.w7(32'h3bc3ac7c),
	.w8(32'h3b5195ab),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be7f9fa),
	.w1(32'h3bae0d44),
	.w2(32'h3abba34b),
	.w3(32'h3b253ada),
	.w4(32'hbc7aa90f),
	.w5(32'hbb62ce1c),
	.w6(32'hbaf94c54),
	.w7(32'h3b196ed9),
	.w8(32'h3b821fd9),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c22e524),
	.w1(32'h3c208371),
	.w2(32'h3cbcdf52),
	.w3(32'h3a3d9042),
	.w4(32'h3ca36a4d),
	.w5(32'h3c3f1128),
	.w6(32'h3c84deaf),
	.w7(32'h3ae3a72d),
	.w8(32'h3bef515d),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd9888d),
	.w1(32'h3bb10b00),
	.w2(32'hbc990776),
	.w3(32'hbc1f4442),
	.w4(32'h3b0b19d3),
	.w5(32'h3c2624a6),
	.w6(32'hbc2c0c29),
	.w7(32'hbc4ce8d9),
	.w8(32'h3c308a00),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb80636e),
	.w1(32'h3cb1a21a),
	.w2(32'h3c054fec),
	.w3(32'hbc46384e),
	.w4(32'h3bb93c33),
	.w5(32'hbc46ac5a),
	.w6(32'h3c12f1ac),
	.w7(32'hbc192412),
	.w8(32'h3b67f156),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8309b8),
	.w1(32'h3b805066),
	.w2(32'h3b3df274),
	.w3(32'h3ab17347),
	.w4(32'h3c5f01c8),
	.w5(32'h3c1f4956),
	.w6(32'h3bdd2265),
	.w7(32'h3cd9f372),
	.w8(32'hba9b76a2),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc08117d),
	.w1(32'h3b72ac66),
	.w2(32'hbc82f147),
	.w3(32'h3c5444c4),
	.w4(32'h3c04b473),
	.w5(32'h3d920437),
	.w6(32'hbc75f944),
	.w7(32'hbc5356dc),
	.w8(32'hbc50f485),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be89a46),
	.w1(32'hbbb6e72f),
	.w2(32'hbcd07f2a),
	.w3(32'h3b44ed10),
	.w4(32'h3b9bc98e),
	.w5(32'hb99dd523),
	.w6(32'hbca23823),
	.w7(32'h3ca332b8),
	.w8(32'h3b316a31),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb1ab5b),
	.w1(32'h3a940953),
	.w2(32'hbbfddcd6),
	.w3(32'hbc936ca6),
	.w4(32'h3d27f747),
	.w5(32'h3b745e1f),
	.w6(32'hbc946197),
	.w7(32'h3b48b018),
	.w8(32'hbbc1cd02),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd083138),
	.w1(32'h3cb89e05),
	.w2(32'h3c390cc0),
	.w3(32'h3d0c8af4),
	.w4(32'hbca484ca),
	.w5(32'hbcc178c6),
	.w6(32'h3b42c059),
	.w7(32'h3c586e5d),
	.w8(32'hbb847eb7),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc316de6),
	.w1(32'hbb3851ab),
	.w2(32'hbac5a794),
	.w3(32'h3cbc0fc3),
	.w4(32'hbc00ab91),
	.w5(32'hbcbe8c81),
	.w6(32'h3a99fd40),
	.w7(32'h3c7c319c),
	.w8(32'hbaa673e1),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1fa0e3),
	.w1(32'hbcdd6e79),
	.w2(32'h3ce34499),
	.w3(32'hbaf3a306),
	.w4(32'h3c7195b5),
	.w5(32'hbb3fe681),
	.w6(32'hbb7563ba),
	.w7(32'h3c08868b),
	.w8(32'h3b94d408),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcd1a7d),
	.w1(32'hbca44b6f),
	.w2(32'h3c8547d6),
	.w3(32'hbba2a932),
	.w4(32'h3cc4a07a),
	.w5(32'h3c99b57e),
	.w6(32'h3bf736ed),
	.w7(32'h3b59b3ae),
	.w8(32'hbcef7e3e),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcaadf6b),
	.w1(32'h3c214048),
	.w2(32'h3b976802),
	.w3(32'hba3d84ed),
	.w4(32'h3c2e3b1c),
	.w5(32'hbca4e753),
	.w6(32'h3aefddff),
	.w7(32'h3c70b6ef),
	.w8(32'h3d3bb475),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b45ad8d),
	.w1(32'hbbd72587),
	.w2(32'h3c7e506a),
	.w3(32'hbbe70e3f),
	.w4(32'h3bd06015),
	.w5(32'h3c432250),
	.w6(32'hbbc80998),
	.w7(32'hbb756176),
	.w8(32'h3c30f5c6),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf64a41),
	.w1(32'h3ba98b9f),
	.w2(32'h3d229245),
	.w3(32'hbc49ff1f),
	.w4(32'h3baf6ec1),
	.w5(32'h3b4ed6fd),
	.w6(32'hbcc5961b),
	.w7(32'hbc9ff76a),
	.w8(32'hbccb01ab),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b42d1c7),
	.w1(32'hbc8743e8),
	.w2(32'h3c162dbf),
	.w3(32'h3c275528),
	.w4(32'h3ba2a289),
	.w5(32'h3b38a284),
	.w6(32'hbbbee198),
	.w7(32'hbadac886),
	.w8(32'h3cc4c422),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98b6e5e),
	.w1(32'hbc81cfdd),
	.w2(32'hbbf679ae),
	.w3(32'hbb92b36b),
	.w4(32'hbc774091),
	.w5(32'h3ba7a519),
	.w6(32'hbbedf022),
	.w7(32'hbcef189c),
	.w8(32'hbbc4a4f3),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c019da8),
	.w1(32'hbc38696a),
	.w2(32'h3c26e01f),
	.w3(32'hbbbcb982),
	.w4(32'hbd099ab2),
	.w5(32'hbc8e6238),
	.w6(32'hbc38ff99),
	.w7(32'hb9c2758c),
	.w8(32'hbb965b14),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8b54dd),
	.w1(32'hbcb5de1d),
	.w2(32'hbc69edba),
	.w3(32'hbbff11f4),
	.w4(32'h3b0e5923),
	.w5(32'h38c2f16a),
	.w6(32'h3c22b66d),
	.w7(32'hbc690d05),
	.w8(32'h3c65899e),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb986f6c),
	.w1(32'hbbdad151),
	.w2(32'h3c8dd0fd),
	.w3(32'h3c6fbebf),
	.w4(32'h394440ed),
	.w5(32'h3c97d91b),
	.w6(32'h3c0c96fb),
	.w7(32'hbc1cac56),
	.w8(32'h3b0b1705),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbece859),
	.w1(32'h398b00a6),
	.w2(32'h3a44376f),
	.w3(32'hbc00cee1),
	.w4(32'h3be4f0ef),
	.w5(32'h3935ab93),
	.w6(32'h39b320b2),
	.w7(32'hbc9a759e),
	.w8(32'h3b06c185),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule