module layer_10_featuremap_479(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7dc2845),
	.w1(32'hb784a1b8),
	.w2(32'hb79e6425),
	.w3(32'hb804cfd2),
	.w4(32'hb8170bf8),
	.w5(32'hb736e631),
	.w6(32'hb7d5db7d),
	.w7(32'hb815d5ea),
	.w8(32'hb6dde27d),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb892970),
	.w1(32'hbbb76bbf),
	.w2(32'hbb8cc48e),
	.w3(32'hbad702d1),
	.w4(32'hbab936a3),
	.w5(32'hbaeef346),
	.w6(32'h3a284588),
	.w7(32'h3a7cd2cf),
	.w8(32'hba00678a),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7b7c4d6),
	.w1(32'hb78c11b2),
	.w2(32'hb7a5603d),
	.w3(32'hb629eb2f),
	.w4(32'h35004c85),
	.w5(32'hb6af5921),
	.w6(32'hb62e8d40),
	.w7(32'h3566c29b),
	.w8(32'hb7142bdb),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba656359),
	.w1(32'hbab5b1cf),
	.w2(32'hbaa00318),
	.w3(32'h38ccd962),
	.w4(32'hba55da0e),
	.w5(32'hb7b63b15),
	.w6(32'h3a3c1540),
	.w7(32'hba19036d),
	.w8(32'hb9e69c53),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba258956),
	.w1(32'hba219d30),
	.w2(32'hb9bbcd7c),
	.w3(32'hba56a330),
	.w4(32'hba436981),
	.w5(32'hb9e20172),
	.w6(32'hba480ab5),
	.w7(32'hba2196c1),
	.w8(32'hb9c69cbd),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h349222a0),
	.w1(32'h378f8b37),
	.w2(32'h37ae5b1f),
	.w3(32'hb6d1be54),
	.w4(32'hb783ebea),
	.w5(32'hb6fc4051),
	.w6(32'hb737bee8),
	.w7(32'hb4b18387),
	.w8(32'h375f43b2),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb12a94b),
	.w1(32'h3aace6c1),
	.w2(32'hb937e1c3),
	.w3(32'h3a8d3634),
	.w4(32'h39b4d425),
	.w5(32'h3b49fd00),
	.w6(32'hbaf2288f),
	.w7(32'h3adc4d9d),
	.w8(32'h3bbe6a24),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8f303f),
	.w1(32'h3c07c357),
	.w2(32'h3bfbb49b),
	.w3(32'hbb264569),
	.w4(32'h3b5bc2e8),
	.w5(32'h3c08ca91),
	.w6(32'hba6f9882),
	.w7(32'hb9ee9442),
	.w8(32'hbb81abc5),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a99ee79),
	.w1(32'hba1e5368),
	.w2(32'h388c70f3),
	.w3(32'hb953dae4),
	.w4(32'hbafdebda),
	.w5(32'hba8193ea),
	.w6(32'hba798666),
	.w7(32'hbae4ea28),
	.w8(32'hba40d84b),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c16b416),
	.w1(32'h3c023e0f),
	.w2(32'h3bc14c29),
	.w3(32'h3b5e87c5),
	.w4(32'h3b43562c),
	.w5(32'h3b65cc7c),
	.w6(32'hbb10f130),
	.w7(32'hbb88a288),
	.w8(32'h3a27d469),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a278fce),
	.w1(32'h3804a9c3),
	.w2(32'h3989a4dc),
	.w3(32'h3a7785e1),
	.w4(32'h36e5e376),
	.w5(32'h3a386575),
	.w6(32'h39756b1b),
	.w7(32'hb9570342),
	.w8(32'h3a0d8162),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3fb963),
	.w1(32'h3b336680),
	.w2(32'h3b1d3f85),
	.w3(32'hbb2b676d),
	.w4(32'hbb18e918),
	.w5(32'hba5279c6),
	.w6(32'hbba78215),
	.w7(32'hbb050eaa),
	.w8(32'h3a8216c5),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c382176),
	.w1(32'h3c3442f9),
	.w2(32'h3bad9602),
	.w3(32'h3bad6b7e),
	.w4(32'h3bdd6745),
	.w5(32'h3bfa55a5),
	.w6(32'hba2c2b0e),
	.w7(32'hb9483818),
	.w8(32'h3b89a8ad),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0d6c6a),
	.w1(32'h39e47ac9),
	.w2(32'hba5172c7),
	.w3(32'hb9ffa9df),
	.w4(32'h3a8c9213),
	.w5(32'h3b3ab0e0),
	.w6(32'hba269243),
	.w7(32'h3aaed2d6),
	.w8(32'h3ab7433a),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af7c8e5),
	.w1(32'hbae9404d),
	.w2(32'hba3e09ea),
	.w3(32'h3a22f35f),
	.w4(32'hbb3b13a9),
	.w5(32'hbb3318f5),
	.w6(32'h3ac922ee),
	.w7(32'hbb332522),
	.w8(32'hbbae238d),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0e69bb),
	.w1(32'h3b4562f3),
	.w2(32'h3a49e3f6),
	.w3(32'h3a86b085),
	.w4(32'h3aa5bba6),
	.w5(32'h3ad75e96),
	.w6(32'hbb82f7c0),
	.w7(32'hbb7ae56c),
	.w8(32'hb980d3e5),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab7f383),
	.w1(32'hba8580b7),
	.w2(32'hba2ee69d),
	.w3(32'hba2a4e1b),
	.w4(32'hba28ba0f),
	.w5(32'hb892a714),
	.w6(32'hb922934f),
	.w7(32'hba117483),
	.w8(32'hba1a340b),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1bfe2a),
	.w1(32'h3be06819),
	.w2(32'hbaabf82e),
	.w3(32'hbba9fac3),
	.w4(32'h3b436b1a),
	.w5(32'h3b110838),
	.w6(32'hbc24c5cc),
	.w7(32'hbbd38793),
	.w8(32'hba81183d),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b92c441),
	.w1(32'h3be69f4a),
	.w2(32'h3b88f5ca),
	.w3(32'h3975cfb4),
	.w4(32'h3bbd57af),
	.w5(32'h3bb2cf88),
	.w6(32'hbb49ebeb),
	.w7(32'hb926a21a),
	.w8(32'h3b693740),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb847c006),
	.w1(32'hb83dbe5d),
	.w2(32'h38d0b1bf),
	.w3(32'h38d0f2e5),
	.w4(32'hb8d5f745),
	.w5(32'h360c8996),
	.w6(32'hb8c9b30c),
	.w7(32'hb93a431e),
	.w8(32'hb90635ea),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb71a7171),
	.w1(32'h38fb6b67),
	.w2(32'h39157160),
	.w3(32'hb7dae0f7),
	.w4(32'hb7d3d2cd),
	.w5(32'h38c01dca),
	.w6(32'hb94ec675),
	.w7(32'h382cef31),
	.w8(32'hb8fb39cf),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb886bdc),
	.w1(32'hbb5e6639),
	.w2(32'hbb26f939),
	.w3(32'hbaab9178),
	.w4(32'hba4a02f4),
	.w5(32'hba9ff99d),
	.w6(32'h3a662006),
	.w7(32'h3a84f973),
	.w8(32'hb9acdb3b),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5bef60),
	.w1(32'h3af03ace),
	.w2(32'h3b6dea50),
	.w3(32'h38418da0),
	.w4(32'hbbc0ed65),
	.w5(32'hbbb4c7e1),
	.w6(32'hbc223a2b),
	.w7(32'hbc3acabc),
	.w8(32'hbb88a7d3),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b79f5bb),
	.w1(32'h3ae14a4f),
	.w2(32'h3acd2cde),
	.w3(32'hbac7ef96),
	.w4(32'hbb56f8ce),
	.w5(32'h374002af),
	.w6(32'hbb740ab9),
	.w7(32'hbbc5319e),
	.w8(32'hbb69b132),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0bc50c),
	.w1(32'hbc138ecb),
	.w2(32'hbbc1f7e0),
	.w3(32'h3b34e435),
	.w4(32'hbb06a901),
	.w5(32'hbb702f67),
	.w6(32'h3c149767),
	.w7(32'h3b860881),
	.w8(32'hba14e5dc),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0e4493),
	.w1(32'hba868f25),
	.w2(32'hbaa102bc),
	.w3(32'h39faae4d),
	.w4(32'hba29c5a8),
	.w5(32'hba1dc0fe),
	.w6(32'h39f8edab),
	.w7(32'hb9d9206c),
	.w8(32'hb8a050a6),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb952e2fb),
	.w1(32'hb9021f29),
	.w2(32'hb94a09f0),
	.w3(32'hb87f987d),
	.w4(32'hb7d01991),
	.w5(32'hb92d17aa),
	.w6(32'hb88ec127),
	.w7(32'hb6e039c1),
	.w8(32'hb8cf0b29),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b39d70c),
	.w1(32'h3b052d0d),
	.w2(32'hbb49c8fc),
	.w3(32'h3b369179),
	.w4(32'h3c7b67f8),
	.w5(32'h3b8eb21b),
	.w6(32'h3b06c0c7),
	.w7(32'h3c2663ae),
	.w8(32'h3bc793d4),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb621ea7),
	.w1(32'hbb2b2137),
	.w2(32'hbadeed90),
	.w3(32'hbb28c353),
	.w4(32'hbb127f1e),
	.w5(32'hbabaf6f7),
	.w6(32'hba9e1a08),
	.w7(32'hbaa5e0e1),
	.w8(32'hbab4c422),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0486ed),
	.w1(32'hbc0a395d),
	.w2(32'hbb85b9e0),
	.w3(32'h3bad58f2),
	.w4(32'h3b807724),
	.w5(32'h3b83d3e4),
	.w6(32'h3b9c705d),
	.w7(32'h3be32f49),
	.w8(32'h3b89ae17),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8820354),
	.w1(32'hb83cae3c),
	.w2(32'hb8456b2c),
	.w3(32'hb84fd803),
	.w4(32'hb847434a),
	.w5(32'hb81f14a5),
	.w6(32'hb8845aa2),
	.w7(32'hb88db1d8),
	.w8(32'hb8805f71),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88ba441),
	.w1(32'hb8b36162),
	.w2(32'hb9593016),
	.w3(32'hb88da70a),
	.w4(32'hb92a6d45),
	.w5(32'hb982c536),
	.w6(32'hb931b063),
	.w7(32'hb99d76cf),
	.w8(32'hb9ada851),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390be54f),
	.w1(32'h394324c1),
	.w2(32'h39febf2d),
	.w3(32'hbb107cc0),
	.w4(32'hbb1ed420),
	.w5(32'hba47ee24),
	.w6(32'hbb8f73ff),
	.w7(32'hbba461da),
	.w8(32'hbb32818a),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a72ab4d),
	.w1(32'hbb03cb82),
	.w2(32'hba440a26),
	.w3(32'h3ae17166),
	.w4(32'h38989b3f),
	.w5(32'hb9eb365a),
	.w6(32'h3b53919c),
	.w7(32'h3a8f8e03),
	.w8(32'h39822c5b),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3bb094),
	.w1(32'h3a239770),
	.w2(32'hb9ab0f32),
	.w3(32'h3a0dc197),
	.w4(32'h3a9ad163),
	.w5(32'h3990ed9a),
	.w6(32'h39b5bf1b),
	.w7(32'h3a143a44),
	.w8(32'h39a28036),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac580f6),
	.w1(32'h3ab3e8af),
	.w2(32'h3aafd221),
	.w3(32'hba3a9933),
	.w4(32'hba6aee6f),
	.w5(32'h3b302f7f),
	.w6(32'hba99e923),
	.w7(32'hbace55a5),
	.w8(32'h3abdeb35),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h356eac80),
	.w1(32'h3b8b3a6b),
	.w2(32'h3bd046b2),
	.w3(32'hba2cbcf7),
	.w4(32'hbc03ae4f),
	.w5(32'hbc1c6a01),
	.w6(32'hba10da0e),
	.w7(32'hbc499b42),
	.w8(32'hbc0a78e7),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4e2d98),
	.w1(32'hbb984e7b),
	.w2(32'hbb92b7ed),
	.w3(32'h3bbf4a23),
	.w4(32'hbb39f744),
	.w5(32'hbc147571),
	.w6(32'h3c3895b5),
	.w7(32'h3ab45071),
	.w8(32'hbc124c51),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb002137),
	.w1(32'hbb13e069),
	.w2(32'hbc1a940c),
	.w3(32'h3b1918a7),
	.w4(32'h3baf8982),
	.w5(32'hbb0ca9ff),
	.w6(32'h3b613711),
	.w7(32'h3bf37543),
	.w8(32'h3b2ec953),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1131de),
	.w1(32'hbb1631c6),
	.w2(32'hba0cd770),
	.w3(32'h39e200b4),
	.w4(32'hb9ffe073),
	.w5(32'h39a65c9c),
	.w6(32'h3ab14927),
	.w7(32'h3a1a003c),
	.w8(32'h39a8bd98),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392c462d),
	.w1(32'h39724a72),
	.w2(32'h391295f7),
	.w3(32'h393fb76c),
	.w4(32'h395543aa),
	.w5(32'h392200b7),
	.w6(32'h383abe22),
	.w7(32'h3915b477),
	.w8(32'h38fccd54),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb68a923b),
	.w1(32'hb62bd6f6),
	.w2(32'hb9228eb3),
	.w3(32'h389c4b72),
	.w4(32'h3710a93b),
	.w5(32'hb94c720b),
	.w6(32'h38c2dfd8),
	.w7(32'h390e73e4),
	.w8(32'hb8dd3d7b),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab93d83),
	.w1(32'h39b05b9a),
	.w2(32'hbb1096f9),
	.w3(32'h3a62331b),
	.w4(32'hbaa2448f),
	.w5(32'hbb093b4e),
	.w6(32'hba11558d),
	.w7(32'hbb043473),
	.w8(32'hbabafa68),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c994186),
	.w1(32'h3c0c60a0),
	.w2(32'h3b66f98c),
	.w3(32'h3ae7bbc5),
	.w4(32'h3b3effe0),
	.w5(32'h3b568886),
	.w6(32'hbc08cba5),
	.w7(32'hbb2399c0),
	.w8(32'h3a80f67e),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba6e5b3),
	.w1(32'hbabfea8a),
	.w2(32'h3906ba84),
	.w3(32'h3b056195),
	.w4(32'hbb4b3030),
	.w5(32'hbadf66aa),
	.w6(32'h3a2ede8d),
	.w7(32'hbba2160e),
	.w8(32'hbb980e12),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9ce7b4),
	.w1(32'h3a94f1c0),
	.w2(32'h3b284e4e),
	.w3(32'hb9b43ef0),
	.w4(32'hbb8006c6),
	.w5(32'h3984faeb),
	.w6(32'hba9d3a83),
	.w7(32'hbbea261e),
	.w8(32'hbbc95549),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3f7447),
	.w1(32'h3ac418ef),
	.w2(32'hba159087),
	.w3(32'h3adfa20f),
	.w4(32'h3a5143a6),
	.w5(32'hba28c404),
	.w6(32'hbaa864c3),
	.w7(32'hbb17281f),
	.w8(32'hbb256607),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc94050),
	.w1(32'h3c577dbf),
	.w2(32'h3bb4a36b),
	.w3(32'hbb0ee8dc),
	.w4(32'h3be8ed8d),
	.w5(32'h3c020731),
	.w6(32'hbc3fce94),
	.w7(32'hbb6897b2),
	.w8(32'h3b573499),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0ff303),
	.w1(32'hb9d4a3c4),
	.w2(32'hb9cc8aa1),
	.w3(32'hb9154c26),
	.w4(32'hb99cad29),
	.w5(32'hb9f73533),
	.w6(32'hb75b5d64),
	.w7(32'hb7872407),
	.w8(32'hb8b5ee84),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b17f7e8),
	.w1(32'h3a87d228),
	.w2(32'h3aab1460),
	.w3(32'h3b006af9),
	.w4(32'h3ac0fb55),
	.w5(32'h3b01da3b),
	.w6(32'h3ae04da5),
	.w7(32'h3abd2551),
	.w8(32'h3b0bdb09),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ba33d9),
	.w1(32'hba17685d),
	.w2(32'h38d9f40f),
	.w3(32'hb98cb5b0),
	.w4(32'hb9ed412e),
	.w5(32'h39ded94d),
	.w6(32'hb9d9f822),
	.w7(32'hb981b7e3),
	.w8(32'h3a0b978c),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bca1d31),
	.w1(32'h3b018aff),
	.w2(32'h3a818622),
	.w3(32'h3aabded1),
	.w4(32'h3a818622),
	.w5(32'h3a48d827),
	.w6(32'h39690988),
	.w7(32'h39ee35b8),
	.w8(32'h3996310d),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a04a25a),
	.w1(32'h3a8021b8),
	.w2(32'h3aa8bdc7),
	.w3(32'hb9e414df),
	.w4(32'hba0135ff),
	.w5(32'h39c01141),
	.w6(32'hba86e7d7),
	.w7(32'hb9b78f86),
	.w8(32'hb9d3f734),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c71ef1e),
	.w1(32'h3c601a51),
	.w2(32'h3b97fa98),
	.w3(32'h3bc16f48),
	.w4(32'h3c06d05e),
	.w5(32'h3b2d600b),
	.w6(32'hbbe84a49),
	.w7(32'hbbc3265d),
	.w8(32'hbaccda9a),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3a2ec9),
	.w1(32'h3b043c51),
	.w2(32'h38050bd7),
	.w3(32'hb8061f7d),
	.w4(32'h3a569cf9),
	.w5(32'h39fbf9fc),
	.w6(32'hb89bb722),
	.w7(32'hba230ed8),
	.w8(32'hba468750),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9421da4),
	.w1(32'hba337a80),
	.w2(32'hb99b0475),
	.w3(32'h38cbc63c),
	.w4(32'hb90413d3),
	.w5(32'hb843002f),
	.w6(32'h39a6dc9e),
	.w7(32'h39acc493),
	.w8(32'h399cd009),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb881a22f),
	.w1(32'hb78b4170),
	.w2(32'hb733f33a),
	.w3(32'hb8496e70),
	.w4(32'hb5d0732f),
	.w5(32'hb82388af),
	.w6(32'hb7a95d01),
	.w7(32'h3788366a),
	.w8(32'hb7c8c340),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38148d3c),
	.w1(32'hb90f03fb),
	.w2(32'hb9bf1f38),
	.w3(32'h39b29d71),
	.w4(32'h3a5145b4),
	.w5(32'hb817e016),
	.w6(32'h39e6cf05),
	.w7(32'h3a3b1244),
	.w8(32'hb800cfdc),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaef1e25),
	.w1(32'hbae99dd9),
	.w2(32'hbabd3407),
	.w3(32'hba8e8b72),
	.w4(32'hba9e26e5),
	.w5(32'hba8f62c9),
	.w6(32'hba2d450e),
	.w7(32'hba6a44cd),
	.w8(32'hba90753f),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9945f7d),
	.w1(32'hb9c653e8),
	.w2(32'hba90fc3c),
	.w3(32'hba0c55c8),
	.w4(32'h390e9a98),
	.w5(32'hb9380be8),
	.w6(32'hb9a14917),
	.w7(32'hb999af8a),
	.w8(32'hb9f65f91),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbad31a),
	.w1(32'h3b2d020b),
	.w2(32'h3a9ba4fb),
	.w3(32'h3a6a18e9),
	.w4(32'h3a4f819f),
	.w5(32'h3a98a15a),
	.w6(32'hbb022f1a),
	.w7(32'hba89d083),
	.w8(32'h399394e6),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2e2733),
	.w1(32'h3ae396a0),
	.w2(32'hbb8952e9),
	.w3(32'h3b087221),
	.w4(32'h3b58ad13),
	.w5(32'hbb01bca6),
	.w6(32'h3b391fe8),
	.w7(32'h3b86a120),
	.w8(32'h3a96261f),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38bb6edc),
	.w1(32'h3810ac56),
	.w2(32'hb703e3ff),
	.w3(32'h38ba3500),
	.w4(32'h388817a1),
	.w5(32'h3569ba7b),
	.w6(32'h3802986f),
	.w7(32'h37247021),
	.w8(32'hb850c25e),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37bbe811),
	.w1(32'h37eda9de),
	.w2(32'h360cf465),
	.w3(32'h383ae4fb),
	.w4(32'h383b5f80),
	.w5(32'h37bec5b8),
	.w6(32'h37d261fa),
	.w7(32'h379f9b77),
	.w8(32'hb76cc8cf),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1a3e9e),
	.w1(32'hb9a39de9),
	.w2(32'hb9250309),
	.w3(32'hb9ff0bad),
	.w4(32'hb98637d3),
	.w5(32'hb852e9a6),
	.w6(32'hb9d1e09d),
	.w7(32'hb97e0c4d),
	.w8(32'hb8f4d096),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb875f8b5),
	.w1(32'hb6edea43),
	.w2(32'hb88da470),
	.w3(32'hb7314de6),
	.w4(32'h37b51bb3),
	.w5(32'hb88068cb),
	.w6(32'hb811832b),
	.w7(32'hb78a1996),
	.w8(32'hb8b04fb3),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c31f358),
	.w1(32'h3c804b32),
	.w2(32'h3a8fc31d),
	.w3(32'h3b196f2e),
	.w4(32'h3c00de6d),
	.w5(32'hbb214317),
	.w6(32'hbbaf7364),
	.w7(32'h39fc4792),
	.w8(32'h3965523a),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb980f48),
	.w1(32'h3aa98730),
	.w2(32'h3bf26f24),
	.w3(32'hbbba6de7),
	.w4(32'hbb6bbb96),
	.w5(32'h3bd37e6e),
	.w6(32'hbc080064),
	.w7(32'hbbd2fc2a),
	.w8(32'hbba3d7b5),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be3009f),
	.w1(32'h3b28ecb4),
	.w2(32'hbb612ca5),
	.w3(32'hbb5e4e6f),
	.w4(32'hbb3f2a0f),
	.w5(32'hbb94ef81),
	.w6(32'hbb85bc59),
	.w7(32'hbaba9ecb),
	.w8(32'hbba81787),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad2fa63),
	.w1(32'hbb564c97),
	.w2(32'hbc03d9bb),
	.w3(32'h3b974618),
	.w4(32'hbbddf640),
	.w5(32'hbc6003ef),
	.w6(32'h3c309ecd),
	.w7(32'h3ae65f43),
	.w8(32'hbbf812bd),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4c92c3),
	.w1(32'h3b8ee316),
	.w2(32'hb89662ff),
	.w3(32'hbb7d797c),
	.w4(32'hbb6ba47a),
	.w5(32'hbbd3d2b1),
	.w6(32'hbb852780),
	.w7(32'h3b6de80d),
	.w8(32'h3b128f8f),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0c21ba),
	.w1(32'hbb8657eb),
	.w2(32'hbbd0bef4),
	.w3(32'hbb88e799),
	.w4(32'hbbe86167),
	.w5(32'hbbc2f166),
	.w6(32'h3aea44ec),
	.w7(32'h3af1e922),
	.w8(32'hbb8d106a),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb11a310),
	.w1(32'h3ae5e8bf),
	.w2(32'hbb97de8d),
	.w3(32'hbbf9c2ea),
	.w4(32'hbad95a24),
	.w5(32'h3a7a724c),
	.w6(32'hbb8409ef),
	.w7(32'hbb149928),
	.w8(32'hbb08e751),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b506c4a),
	.w1(32'h3a714b34),
	.w2(32'h3b625320),
	.w3(32'hba20b9b1),
	.w4(32'h3ba9bac1),
	.w5(32'h3c1a3857),
	.w6(32'hbba902ef),
	.w7(32'hbb3b5d3d),
	.w8(32'h3a149350),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7741c6),
	.w1(32'h3add7528),
	.w2(32'hba93ab76),
	.w3(32'h3bc20ccf),
	.w4(32'hbbc688c3),
	.w5(32'hbb45b9e1),
	.w6(32'h3bd8a151),
	.w7(32'hb9c545b5),
	.w8(32'hbb071b03),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b969fcd),
	.w1(32'h3c0deb80),
	.w2(32'h3b743ee9),
	.w3(32'hbac9ee4f),
	.w4(32'h3b3f69b4),
	.w5(32'h3c34ba71),
	.w6(32'h379adc1a),
	.w7(32'hba7b4661),
	.w8(32'hbb58c8ef),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f2fed),
	.w1(32'h3c0eb153),
	.w2(32'h3c2c346e),
	.w3(32'hbb551ac1),
	.w4(32'hba9a1559),
	.w5(32'h3c0d2985),
	.w6(32'hbc10b18e),
	.w7(32'h39369c64),
	.w8(32'h3bec7fe7),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3addb931),
	.w1(32'h3be1331b),
	.w2(32'hbc091ddd),
	.w3(32'h3ba62533),
	.w4(32'h3c239aae),
	.w5(32'h3cc8b788),
	.w6(32'h3bc3c7cb),
	.w7(32'h3b4751a3),
	.w8(32'hbc0a4d59),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcac7b0),
	.w1(32'h3c31998b),
	.w2(32'h396ebba6),
	.w3(32'h3c4df8c9),
	.w4(32'h3bd62eeb),
	.w5(32'h3c129ce7),
	.w6(32'hbabca64e),
	.w7(32'h3abbd749),
	.w8(32'hbc0856ad),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8e3276),
	.w1(32'h3bf53305),
	.w2(32'h39761734),
	.w3(32'h3b8b6b79),
	.w4(32'hbb6ea6ae),
	.w5(32'hbba523a1),
	.w6(32'hbc0f12ec),
	.w7(32'h3b600af5),
	.w8(32'h3b4d0a94),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb1d2ee),
	.w1(32'h3c42d978),
	.w2(32'h3bd026f2),
	.w3(32'h3b61995f),
	.w4(32'h3b867b09),
	.w5(32'h3bb6c818),
	.w6(32'h3b1ad8e1),
	.w7(32'hba77dcda),
	.w8(32'hbb59f464),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1fc982),
	.w1(32'h3b2a9cca),
	.w2(32'h3b1c58cb),
	.w3(32'h3c078051),
	.w4(32'h3b87fa67),
	.w5(32'h396f4580),
	.w6(32'hba74f4ef),
	.w7(32'hbaef41fc),
	.w8(32'h3b16fd41),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a803609),
	.w1(32'hbb8ddf75),
	.w2(32'hbb04e8f7),
	.w3(32'h3b14197b),
	.w4(32'hbb0a9d35),
	.w5(32'hbbcaa89c),
	.w6(32'hbab6790d),
	.w7(32'h3b976a6f),
	.w8(32'h3a215347),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b37859b),
	.w1(32'h3b7fa5a9),
	.w2(32'hb960edc6),
	.w3(32'hbb5fb556),
	.w4(32'hb480a5a8),
	.w5(32'hbbf9eec0),
	.w6(32'h3a33943c),
	.w7(32'h3b5e9d4c),
	.w8(32'h3b8d640f),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b951817),
	.w1(32'h3aad0c97),
	.w2(32'h3b09f9e0),
	.w3(32'hbbaa4108),
	.w4(32'h3b856a06),
	.w5(32'h39b9e7a5),
	.w6(32'h3b816e17),
	.w7(32'h39880e6a),
	.w8(32'h3bd3126b),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf645cd),
	.w1(32'hbbad1585),
	.w2(32'hbb1f9544),
	.w3(32'h3aa6ae6d),
	.w4(32'hbbb3be9f),
	.w5(32'hbbae0e2f),
	.w6(32'h3a82f814),
	.w7(32'hbbbf0e53),
	.w8(32'h390283ef),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb67ca37),
	.w1(32'h3c003b1a),
	.w2(32'hbac82a94),
	.w3(32'hba8b7c9d),
	.w4(32'h3bc0c8fa),
	.w5(32'h3c8e497f),
	.w6(32'h3aae49a0),
	.w7(32'hbb8ea41f),
	.w8(32'hbbb15b2f),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf761d7),
	.w1(32'hba4f0cc4),
	.w2(32'hbb290bde),
	.w3(32'h3c3bd6e7),
	.w4(32'h3c00a7c8),
	.w5(32'h3cd55377),
	.w6(32'h3b51e074),
	.w7(32'hbbb6d086),
	.w8(32'hbb82cf3d),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbdff05),
	.w1(32'hbbed6db8),
	.w2(32'hba20be6b),
	.w3(32'h3bf24e4a),
	.w4(32'hbbbf62a9),
	.w5(32'h3aaac70c),
	.w6(32'h3b42c6eb),
	.w7(32'hbba182ab),
	.w8(32'hbbaaad7f),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be8af9d),
	.w1(32'h3bddfa2c),
	.w2(32'h3b574ae1),
	.w3(32'hbc19e33f),
	.w4(32'h3b1529ab),
	.w5(32'h3c0ffc6d),
	.w6(32'hbc375949),
	.w7(32'h3a7053f6),
	.w8(32'hb9c05a37),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3f0feb),
	.w1(32'hbb248499),
	.w2(32'hbbbf58b4),
	.w3(32'h3be561e0),
	.w4(32'h3b96ee22),
	.w5(32'hbbaaba96),
	.w6(32'hbb1e1567),
	.w7(32'h3b7458b3),
	.w8(32'h3bad3c2e),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4febd3),
	.w1(32'h3c4bfdb1),
	.w2(32'h3bafc4cc),
	.w3(32'hbb974e51),
	.w4(32'hbc3267af),
	.w5(32'hbc826220),
	.w6(32'hbb58dc6b),
	.w7(32'h3ab63504),
	.w8(32'hbb5659d3),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaab797c),
	.w1(32'hbc57f183),
	.w2(32'hbc4d236e),
	.w3(32'hbbf41de4),
	.w4(32'hbc085c71),
	.w5(32'hbc1838bb),
	.w6(32'h3aeeee34),
	.w7(32'h3b22d06a),
	.w8(32'h3a132f80),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c57fd35),
	.w1(32'h3c7df490),
	.w2(32'h3c45085e),
	.w3(32'hbc4d66d2),
	.w4(32'hbab2d3af),
	.w5(32'hb90b3a76),
	.w6(32'hbc29662e),
	.w7(32'hbb47fac0),
	.w8(32'hbb63e41a),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0b3b8a),
	.w1(32'h3b2a0b3d),
	.w2(32'h3ad985b6),
	.w3(32'hb9fe47b0),
	.w4(32'hbba9365c),
	.w5(32'hbbcc6da8),
	.w6(32'hbc2abeb7),
	.w7(32'hbad2d7bb),
	.w8(32'hba8430ce),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc35ab9),
	.w1(32'hbbe77a08),
	.w2(32'h3a86fbf5),
	.w3(32'h3bb2b356),
	.w4(32'hba87f869),
	.w5(32'hbc4d01ac),
	.w6(32'h3c0e7a9a),
	.w7(32'hbb7a96b3),
	.w8(32'hbb320ebc),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9efac19),
	.w1(32'hbbd2a391),
	.w2(32'h3b421bac),
	.w3(32'hbba199a7),
	.w4(32'h3b4638e6),
	.w5(32'hbc277baf),
	.w6(32'hbb82fd31),
	.w7(32'hbbbea6cb),
	.w8(32'hbbb3aac2),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c323094),
	.w1(32'h3b8e735c),
	.w2(32'h3b1de6c9),
	.w3(32'h3b4bc016),
	.w4(32'h3bb3e85b),
	.w5(32'h3a85a37c),
	.w6(32'hbb113e43),
	.w7(32'h3aaed613),
	.w8(32'hbab23c3b),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1eabd0),
	.w1(32'h3c1fb217),
	.w2(32'h3b931555),
	.w3(32'h391fbaa7),
	.w4(32'hbb3d5ab9),
	.w5(32'hbbbef550),
	.w6(32'hbb94d45d),
	.w7(32'hba95fd03),
	.w8(32'h3a8953bc),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbea50d8),
	.w1(32'hbb178f98),
	.w2(32'h3b030b66),
	.w3(32'hbbd4d212),
	.w4(32'hbc39acb6),
	.w5(32'hbc0ec37d),
	.w6(32'hbb524441),
	.w7(32'hbb9f705c),
	.w8(32'hbb9f8f70),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bed7332),
	.w1(32'hbb1b40dd),
	.w2(32'hbb3e9745),
	.w3(32'h3b97bf5b),
	.w4(32'hbadb276a),
	.w5(32'h3af613cf),
	.w6(32'h3c292ed9),
	.w7(32'hbbb3eef8),
	.w8(32'hbc022295),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8ee01b),
	.w1(32'hbbbd4e6e),
	.w2(32'h3b429211),
	.w3(32'h3c535463),
	.w4(32'hbbb1048d),
	.w5(32'hbbd0aaa7),
	.w6(32'h3c4e665c),
	.w7(32'hbb84d3bc),
	.w8(32'hba639a3e),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd0885f),
	.w1(32'h3c5b3a6a),
	.w2(32'h3b44b005),
	.w3(32'hbb1e74b6),
	.w4(32'hb9f258cd),
	.w5(32'h3b887fcd),
	.w6(32'hbc1063fb),
	.w7(32'hbc3c74ed),
	.w8(32'hbb0f0723),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3add87cb),
	.w1(32'h394e3e0a),
	.w2(32'hbb983650),
	.w3(32'h3baab188),
	.w4(32'hbaa425ef),
	.w5(32'hbbe5fa15),
	.w6(32'h3b013ec8),
	.w7(32'hbacb43c1),
	.w8(32'hbbb94d31),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1ed9c3),
	.w1(32'h3b665c78),
	.w2(32'h3b4d3615),
	.w3(32'h3bbb1be7),
	.w4(32'hbc3fca86),
	.w5(32'hbc62a58d),
	.w6(32'hbba3713a),
	.w7(32'hbb860722),
	.w8(32'hbb794bd6),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a91addf),
	.w1(32'h3a1c8651),
	.w2(32'h3b61625c),
	.w3(32'hbc4470e9),
	.w4(32'hba260110),
	.w5(32'h3a416ae4),
	.w6(32'h3bbbe54f),
	.w7(32'h3b5f5630),
	.w8(32'h3c0aede9),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb65e63a),
	.w1(32'hbb22a409),
	.w2(32'hbb23dfd2),
	.w3(32'hbb25e288),
	.w4(32'hba874dd6),
	.w5(32'hbaaf8a64),
	.w6(32'h3b0049df),
	.w7(32'hbb480851),
	.w8(32'hbb890660),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba900197),
	.w1(32'h3b0c8ef1),
	.w2(32'hba16e446),
	.w3(32'h3ad9735e),
	.w4(32'h3911d987),
	.w5(32'hbb3d45f4),
	.w6(32'hbaa88259),
	.w7(32'h3b2a8ce9),
	.w8(32'h3b73854b),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b87c0ed),
	.w1(32'h39025f9b),
	.w2(32'h39a9c588),
	.w3(32'hbbc4e88b),
	.w4(32'hbb46e776),
	.w5(32'hbaa83f3b),
	.w6(32'hbbd3131b),
	.w7(32'h3b391c41),
	.w8(32'h3b812ac2),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb008510),
	.w1(32'hbb5ddf62),
	.w2(32'hb9b70eb2),
	.w3(32'hbbf8d923),
	.w4(32'hbb20d0f1),
	.w5(32'hba088c92),
	.w6(32'h3b492c85),
	.w7(32'h3c08240e),
	.w8(32'h3c764610),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c050b5c),
	.w1(32'h3c07f0e2),
	.w2(32'h3b69b3f5),
	.w3(32'hbb365b25),
	.w4(32'h3abdd97f),
	.w5(32'hbbb99877),
	.w6(32'h3ba54cfa),
	.w7(32'h3bdc3554),
	.w8(32'h3bb92000),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfd10b2),
	.w1(32'h3a66a811),
	.w2(32'h3b4ca32c),
	.w3(32'h3bb4bbee),
	.w4(32'hbad69ff1),
	.w5(32'hbc0e4675),
	.w6(32'h3c3c4a8c),
	.w7(32'h3b82be2b),
	.w8(32'hbb7549e1),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb010666),
	.w1(32'h3b389020),
	.w2(32'h3bed0e89),
	.w3(32'h3b469db8),
	.w4(32'h3a036113),
	.w5(32'h3bb21684),
	.w6(32'h3b8adbd4),
	.w7(32'hbb6280e5),
	.w8(32'h3af850ef),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8a2801),
	.w1(32'h3c3eaeab),
	.w2(32'h3b6e99e8),
	.w3(32'h3c746c45),
	.w4(32'hbb9427dd),
	.w5(32'hbc004897),
	.w6(32'h3c140d9c),
	.w7(32'hbbab4f25),
	.w8(32'hbb544cff),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c303823),
	.w1(32'h3819defb),
	.w2(32'h3b0173db),
	.w3(32'hbb515f0f),
	.w4(32'hbab81aa7),
	.w5(32'hbb669143),
	.w6(32'h3ac9d5bc),
	.w7(32'hbad072c8),
	.w8(32'hbafeaad4),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfbaf80),
	.w1(32'h3b90cf23),
	.w2(32'h39c24c94),
	.w3(32'hbad27f97),
	.w4(32'hbb3c67f5),
	.w5(32'hbb55ed3e),
	.w6(32'hbb85cfc4),
	.w7(32'h3ad7982a),
	.w8(32'hb90da9ad),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af47dac),
	.w1(32'hbb2a3854),
	.w2(32'h3a3c73b2),
	.w3(32'hba29a11b),
	.w4(32'hba3b689e),
	.w5(32'hbb50337b),
	.w6(32'hb8e04748),
	.w7(32'hba8fce22),
	.w8(32'h3bdbe926),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b307b2a),
	.w1(32'hbbbfb3a2),
	.w2(32'hbaf39b93),
	.w3(32'hbb362b91),
	.w4(32'hbb58e66c),
	.w5(32'hbc2494ad),
	.w6(32'hba948041),
	.w7(32'h3c32e907),
	.w8(32'h3a36cb90),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b562db4),
	.w1(32'hbbdfd3e5),
	.w2(32'hbc24bbdd),
	.w3(32'hbc4937b0),
	.w4(32'hbba257ea),
	.w5(32'h3c885763),
	.w6(32'hbbf239f6),
	.w7(32'hbc004a7a),
	.w8(32'hbbef0885),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc02b04b),
	.w1(32'hb9ef31bd),
	.w2(32'hbb09fc46),
	.w3(32'h3b49089f),
	.w4(32'hbbf4ae17),
	.w5(32'hbc85b789),
	.w6(32'hba0ad655),
	.w7(32'hbbd1cadb),
	.w8(32'hbc1c92ca),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb5c64f),
	.w1(32'h3ac9a65b),
	.w2(32'h3b2ceb17),
	.w3(32'hbb566e8e),
	.w4(32'h3af874d1),
	.w5(32'h3b6cfc7c),
	.w6(32'hbb824b94),
	.w7(32'hbb4c2432),
	.w8(32'h3b74fd24),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0136fe),
	.w1(32'h3bf4cc72),
	.w2(32'h3a86ee0b),
	.w3(32'hb9867830),
	.w4(32'hbb8b3da8),
	.w5(32'hbb15dae0),
	.w6(32'h3a29a421),
	.w7(32'hbbcf5374),
	.w8(32'h3ac1bc3c),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb789512),
	.w1(32'hbb9705bb),
	.w2(32'hbb2d2f33),
	.w3(32'h39e1ec29),
	.w4(32'h3a844f66),
	.w5(32'hbbad56ba),
	.w6(32'h3b441bf4),
	.w7(32'hba803e4d),
	.w8(32'h3aaf4df8),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b582247),
	.w1(32'h3a149067),
	.w2(32'h3c071bad),
	.w3(32'h3bbf7b85),
	.w4(32'hbb55023e),
	.w5(32'hbc04b48d),
	.w6(32'h3b17de8a),
	.w7(32'hba78bcf9),
	.w8(32'h3b53456d),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1efa1f),
	.w1(32'hbb9ff530),
	.w2(32'hba67d4d5),
	.w3(32'h3b6b35ca),
	.w4(32'hba500990),
	.w5(32'hba3d9be6),
	.w6(32'h3bf9d6b3),
	.w7(32'h3be5dc05),
	.w8(32'h3bd7e911),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ab27d4),
	.w1(32'h3a829203),
	.w2(32'hbb881f98),
	.w3(32'hbc017e5b),
	.w4(32'hbc01ac50),
	.w5(32'hbc1130fa),
	.w6(32'h3a9855df),
	.w7(32'h3a8ccf51),
	.w8(32'hbba7018f),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadd2fdf),
	.w1(32'hbbc0bf5d),
	.w2(32'h3ac0f645),
	.w3(32'hbbccd8e3),
	.w4(32'hbbbfc00b),
	.w5(32'hbb691bc9),
	.w6(32'hbb528e74),
	.w7(32'h3b1946fc),
	.w8(32'hbb1eee8e),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb85eafc),
	.w1(32'hbb178c8e),
	.w2(32'h3bc24b12),
	.w3(32'hb9ff0d94),
	.w4(32'hb97cd5c7),
	.w5(32'h3c26f5f7),
	.w6(32'hbba2e68e),
	.w7(32'hbaaac486),
	.w8(32'hbac5ae27),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c446f6c),
	.w1(32'h3c3ed1d1),
	.w2(32'h3bbac899),
	.w3(32'hbb01eea5),
	.w4(32'h3bb1d33f),
	.w5(32'h3bba5973),
	.w6(32'hbc20ca11),
	.w7(32'hba38141a),
	.w8(32'hbb131d37),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e77292),
	.w1(32'h3c04773d),
	.w2(32'h3ac4b899),
	.w3(32'h3af8454a),
	.w4(32'hbadf578c),
	.w5(32'h3a9deb4d),
	.w6(32'hbb1b0040),
	.w7(32'h3af3ad96),
	.w8(32'hbb236c2e),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb82269),
	.w1(32'hbaf97233),
	.w2(32'hbbf15e3c),
	.w3(32'h3bd703e6),
	.w4(32'h3b82a668),
	.w5(32'h3c42a73a),
	.w6(32'h3b4b0466),
	.w7(32'hb9a0f6dc),
	.w8(32'hba643766),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc130d9a),
	.w1(32'h3b49409d),
	.w2(32'hbaf8e4fa),
	.w3(32'hbb97be98),
	.w4(32'hbc308781),
	.w5(32'hbc8304a3),
	.w6(32'hbbf66ab9),
	.w7(32'h3a833745),
	.w8(32'hbc40a7a7),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baa4a86),
	.w1(32'h3abc8f52),
	.w2(32'h3a2eec90),
	.w3(32'hbbb45848),
	.w4(32'hbb4a3dbe),
	.w5(32'hbbbb62a0),
	.w6(32'hbbb3d2a8),
	.w7(32'h3b5736ea),
	.w8(32'hba2220b8),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3947a9d3),
	.w1(32'h3b629129),
	.w2(32'h3c278f6b),
	.w3(32'hb8f40b23),
	.w4(32'hbaaa0c69),
	.w5(32'hbba555b7),
	.w6(32'hba59b99a),
	.w7(32'hbaec53a0),
	.w8(32'hbb945d08),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c61a0e2),
	.w1(32'h3c3da5ae),
	.w2(32'h3bf77507),
	.w3(32'h39f8bd0c),
	.w4(32'h3c91530e),
	.w5(32'h3cf86f96),
	.w6(32'hbbc2cac4),
	.w7(32'hbb8d0667),
	.w8(32'hbae4f1b1),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab5cc63),
	.w1(32'h3c1692de),
	.w2(32'h3bfe8aa4),
	.w3(32'h3ca440ea),
	.w4(32'h3b8519a1),
	.w5(32'h3c02ee8a),
	.w6(32'h3c5a1c4f),
	.w7(32'hba9d8683),
	.w8(32'hbab1e373),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bab7ccb),
	.w1(32'hbb41f215),
	.w2(32'h3a9135e6),
	.w3(32'h3c80bc6f),
	.w4(32'hbc12bba2),
	.w5(32'hbc5b1f06),
	.w6(32'hb99046d3),
	.w7(32'hbc1adae9),
	.w8(32'hbb833e06),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8dad11),
	.w1(32'h3bf71025),
	.w2(32'h3b8dc5cc),
	.w3(32'hbb7e779f),
	.w4(32'h38c955bd),
	.w5(32'hbb09d431),
	.w6(32'hbc0d2005),
	.w7(32'h3b4fd30a),
	.w8(32'h3bf27a48),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3f79c0),
	.w1(32'hbb78aa6e),
	.w2(32'h3b614036),
	.w3(32'hbc05536b),
	.w4(32'hb8cbf4ae),
	.w5(32'h3b7103f6),
	.w6(32'h3b87d8f6),
	.w7(32'h3b0cbe91),
	.w8(32'h3c03a429),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2012a8),
	.w1(32'h3b3198a4),
	.w2(32'h3b8e05a6),
	.w3(32'h3b7e7f7e),
	.w4(32'hbaba432e),
	.w5(32'h39a0ff42),
	.w6(32'h3a7024af),
	.w7(32'hbb7a43ae),
	.w8(32'h3b7ee2aa),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9aefa5c),
	.w1(32'h3b08790d),
	.w2(32'hbb66d359),
	.w3(32'h3b3567e8),
	.w4(32'hbc41f805),
	.w5(32'hbc7375c2),
	.w6(32'h3b6fb8b0),
	.w7(32'hbb8f4b0a),
	.w8(32'hbc1f2e3c),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f61fe),
	.w1(32'hbb87b25c),
	.w2(32'hbbf217cd),
	.w3(32'hbb99748b),
	.w4(32'h3c0cc173),
	.w5(32'h3c0eaa7c),
	.w6(32'hba6efcee),
	.w7(32'hb864719a),
	.w8(32'h3c0b98d6),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4fd883),
	.w1(32'hbb069429),
	.w2(32'h3b8b5833),
	.w3(32'h3acfcf54),
	.w4(32'h3a92e056),
	.w5(32'hbb38b085),
	.w6(32'hba99f6f7),
	.w7(32'h3ae0eff7),
	.w8(32'hbb40fb90),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba7ed0d),
	.w1(32'h3ad79424),
	.w2(32'h39b31fde),
	.w3(32'hbb39a6e1),
	.w4(32'hba8ce7b2),
	.w5(32'hbb64d7c7),
	.w6(32'h3a46e8b8),
	.w7(32'hbae3229b),
	.w8(32'hbb2a861f),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb39e59c),
	.w1(32'h3b497713),
	.w2(32'hba1bdd16),
	.w3(32'hbb418b9d),
	.w4(32'h3afe2ca0),
	.w5(32'h3b637536),
	.w6(32'h3a8d06d3),
	.w7(32'h3af591bc),
	.w8(32'h3af18b8f),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0955e7),
	.w1(32'h3b48e186),
	.w2(32'h3a24ee96),
	.w3(32'h3b9277e4),
	.w4(32'h3b88930b),
	.w5(32'h3b5eb099),
	.w6(32'h3b5ddcf7),
	.w7(32'h399a4e25),
	.w8(32'h38cb4170),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9e598a),
	.w1(32'hbb4b53f8),
	.w2(32'h3b9f97ea),
	.w3(32'h3a2268c8),
	.w4(32'hbbb05020),
	.w5(32'hbc06326b),
	.w6(32'h3aa4e188),
	.w7(32'hbb3f1290),
	.w8(32'h3a138166),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4be160),
	.w1(32'h3bcf0612),
	.w2(32'hbb55c8e5),
	.w3(32'h3af25855),
	.w4(32'h3c22b6bd),
	.w5(32'h3b6f9a63),
	.w6(32'hb8cfce6a),
	.w7(32'h3b978e9e),
	.w8(32'h3bb63fda),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3fa5f2),
	.w1(32'hbb7daf58),
	.w2(32'h3a3a7e50),
	.w3(32'hbc2f24bb),
	.w4(32'hbb863745),
	.w5(32'hbbd2cebd),
	.w6(32'hbb67087a),
	.w7(32'hbba63f80),
	.w8(32'hbbfae0ff),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1512f9),
	.w1(32'h39bfa938),
	.w2(32'h3aec8a2d),
	.w3(32'h38f62ea4),
	.w4(32'h3ad48865),
	.w5(32'hbaa55898),
	.w6(32'hbc0bc14c),
	.w7(32'hbb18d109),
	.w8(32'h3a21f949),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b601332),
	.w1(32'hbb9254c9),
	.w2(32'hba0c85c9),
	.w3(32'h3ae3f633),
	.w4(32'hbbccc13b),
	.w5(32'hbb02e960),
	.w6(32'h3b9a2f2c),
	.w7(32'hbbdd5500),
	.w8(32'h3a122a1f),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb4f5c7),
	.w1(32'h3c3226c6),
	.w2(32'h3bf07e79),
	.w3(32'hbbd1cdad),
	.w4(32'hba696dd6),
	.w5(32'h3acda81a),
	.w6(32'hbc2f6c9b),
	.w7(32'hbae5eb1c),
	.w8(32'h3ac4b0c5),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0aefac),
	.w1(32'h3bda1c18),
	.w2(32'h3b47025d),
	.w3(32'h3b61f825),
	.w4(32'h3be11d71),
	.w5(32'hbbcf1f4e),
	.w6(32'h3c0b9661),
	.w7(32'h3b7d91fc),
	.w8(32'h3b873cd8),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf48283),
	.w1(32'h3bff70d3),
	.w2(32'h3bcc7720),
	.w3(32'h3ad7ab8b),
	.w4(32'h39a0394b),
	.w5(32'h3b2dc15f),
	.w6(32'h3b469c74),
	.w7(32'h3c05cc03),
	.w8(32'h3bb40533),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be36dd8),
	.w1(32'h3a8b3de7),
	.w2(32'h3b5eb270),
	.w3(32'hb88a9334),
	.w4(32'h3c0504a4),
	.w5(32'h3a99562d),
	.w6(32'h3bc64845),
	.w7(32'hbbe7d45c),
	.w8(32'hbbe822ff),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf9ef71),
	.w1(32'h3be8f1e5),
	.w2(32'h3b75b38c),
	.w3(32'h3be441a6),
	.w4(32'h3b71c22e),
	.w5(32'hba0b2f78),
	.w6(32'h3b01f9c7),
	.w7(32'h38ca2e7f),
	.w8(32'h3b140b03),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b471e77),
	.w1(32'hbb811a9f),
	.w2(32'hbb3b3eb3),
	.w3(32'hbacdf91a),
	.w4(32'hbbf2185d),
	.w5(32'hbbe55b51),
	.w6(32'hbb5cc59f),
	.w7(32'hba369d77),
	.w8(32'hbb48d95d),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbad84bd),
	.w1(32'hbbe98cf3),
	.w2(32'hbb92b347),
	.w3(32'hbb5266f3),
	.w4(32'h3acb8d93),
	.w5(32'h3b99c192),
	.w6(32'h3af9b9e1),
	.w7(32'h3aeae812),
	.w8(32'hbb382703),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb36f5cb),
	.w1(32'hbba35e16),
	.w2(32'hbbe05637),
	.w3(32'h3b1fabfa),
	.w4(32'hbb20f386),
	.w5(32'hb8e8ecbd),
	.w6(32'hbbbf4026),
	.w7(32'h3bb320f3),
	.w8(32'hbb2e2685),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb895b27),
	.w1(32'h3be46ed5),
	.w2(32'hbb0eb8a5),
	.w3(32'hbc090c3d),
	.w4(32'h3b949ff5),
	.w5(32'h3bace09a),
	.w6(32'h3a34b24b),
	.w7(32'hbb082bbe),
	.w8(32'hbb82ce40),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8a9545),
	.w1(32'h3c993811),
	.w2(32'h3c4a2266),
	.w3(32'h3bad9ff3),
	.w4(32'h3c488c10),
	.w5(32'h3cad4c27),
	.w6(32'hbb635df5),
	.w7(32'hbb0e15b7),
	.w8(32'hba97d4d5),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3687e3),
	.w1(32'h3be51675),
	.w2(32'h3b988c66),
	.w3(32'h3c96abc7),
	.w4(32'h3a9107b7),
	.w5(32'h3b83e1d9),
	.w6(32'h3a6d66d8),
	.w7(32'h3b8475e2),
	.w8(32'h3b974b4d),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6c7809),
	.w1(32'hbbc800bb),
	.w2(32'hbbe365cb),
	.w3(32'h3c3e095b),
	.w4(32'h3b29b3c5),
	.w5(32'hbba7177d),
	.w6(32'h3c2f09da),
	.w7(32'h3b924e6f),
	.w8(32'h3b2ba29d),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6bd487),
	.w1(32'h3b6b2476),
	.w2(32'hbab1900a),
	.w3(32'hbb58d0d6),
	.w4(32'hbaa224d2),
	.w5(32'hba87659a),
	.w6(32'hba553a4d),
	.w7(32'h3b4e73ba),
	.w8(32'h391ee30e),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3cc356),
	.w1(32'hbb7b31aa),
	.w2(32'h3ac80004),
	.w3(32'hbbcc3f4a),
	.w4(32'h3b96de29),
	.w5(32'h3bf4f35b),
	.w6(32'hbb89924f),
	.w7(32'h3b4fc876),
	.w8(32'h3aadbcd3),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acb9c4e),
	.w1(32'h3b95071c),
	.w2(32'hbba4595d),
	.w3(32'h3b0944e5),
	.w4(32'hb8be6cd6),
	.w5(32'h3c336a1c),
	.w6(32'h3b9c4bc2),
	.w7(32'hbbcb893c),
	.w8(32'hbbc156ee),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6a63f3),
	.w1(32'hbb6af5ea),
	.w2(32'h3aaf01c2),
	.w3(32'h3c4848ec),
	.w4(32'hbbb7a193),
	.w5(32'hbb5fa63c),
	.w6(32'h38387c9b),
	.w7(32'hbbc24624),
	.w8(32'h3c182a39),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9af27a),
	.w1(32'h3bfc000f),
	.w2(32'hbb110da3),
	.w3(32'hbb9c20ff),
	.w4(32'h3ad5e50f),
	.w5(32'h3812d314),
	.w6(32'hb9583614),
	.w7(32'hbb9c69a7),
	.w8(32'hbbe5cb5d),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b698442),
	.w1(32'h3b7e0973),
	.w2(32'h3c020b53),
	.w3(32'h3b9209a8),
	.w4(32'hbb82c8bb),
	.w5(32'hbb48e75e),
	.w6(32'hbb15280a),
	.w7(32'hbbd8414a),
	.w8(32'hbc0a6c53),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2ac006),
	.w1(32'hbc12380b),
	.w2(32'hbb069cb8),
	.w3(32'hbb977c08),
	.w4(32'hbb8206ec),
	.w5(32'hbc81ab9b),
	.w6(32'hbba700d1),
	.w7(32'hbbd0911b),
	.w8(32'hbbc0b7b9),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba41fbb1),
	.w1(32'hb936f1ee),
	.w2(32'hbb0961a6),
	.w3(32'hbb6c19de),
	.w4(32'hbbfbb66c),
	.w5(32'hbc3653d0),
	.w6(32'hbb5afd61),
	.w7(32'hba4ecf7f),
	.w8(32'hbbef817e),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb28a2b8),
	.w1(32'h3c1538ac),
	.w2(32'h3bb174ba),
	.w3(32'hbc222ccb),
	.w4(32'h3b5a5648),
	.w5(32'hb980178f),
	.w6(32'hbc0abebd),
	.w7(32'hbb1a9c22),
	.w8(32'hba0712d7),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca3e37f),
	.w1(32'h3c63ae0f),
	.w2(32'h3a97d01b),
	.w3(32'hbac9575b),
	.w4(32'h3b3c4f4a),
	.w5(32'hbbeef260),
	.w6(32'hbb8a8923),
	.w7(32'hbacecae0),
	.w8(32'h3ae865a5),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0b6ee9),
	.w1(32'h3b7265e4),
	.w2(32'h3a94e196),
	.w3(32'h3a96f293),
	.w4(32'h3aba0d2a),
	.w5(32'h3a968202),
	.w6(32'hbb7efb8a),
	.w7(32'hbaa4fcca),
	.w8(32'h38b8acb9),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcf5c21),
	.w1(32'hbb2ea7aa),
	.w2(32'h3a1f2cf7),
	.w3(32'hbb13c1f8),
	.w4(32'hbb87056f),
	.w5(32'hba3f43ae),
	.w6(32'hbaee650e),
	.w7(32'hbb3325a6),
	.w8(32'h3a6b8f2d),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acc8dbd),
	.w1(32'hbb78a5e2),
	.w2(32'hbb06c9e4),
	.w3(32'hbbc518f7),
	.w4(32'hbb9c0150),
	.w5(32'hbbf539d5),
	.w6(32'hbbbff5ea),
	.w7(32'hbb76f42f),
	.w8(32'hbaf9d01b),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8b8d53),
	.w1(32'h3b3ec3d2),
	.w2(32'h3b9ebf0d),
	.w3(32'hba926e65),
	.w4(32'h3b5dbae8),
	.w5(32'h39a7ab6c),
	.w6(32'hbb8f9fc1),
	.w7(32'hba5ad8f3),
	.w8(32'h3a05ae36),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b91f7df),
	.w1(32'h3bb4ef9b),
	.w2(32'h3b77c56c),
	.w3(32'h3b4091a1),
	.w4(32'h3b8d54fe),
	.w5(32'h3b0bed13),
	.w6(32'hb8c5582e),
	.w7(32'h3916fd61),
	.w8(32'hbac41e73),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf67b00),
	.w1(32'hba26de76),
	.w2(32'h3a7ebd0b),
	.w3(32'h3b2f21e6),
	.w4(32'hbb5e55e9),
	.w5(32'hbbc63330),
	.w6(32'h3b232f25),
	.w7(32'h3bf73cb2),
	.w8(32'h3a6ac946),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39626be5),
	.w1(32'hbbc613f5),
	.w2(32'hbb965862),
	.w3(32'hb952996c),
	.w4(32'hbaea6c35),
	.w5(32'hbb80139c),
	.w6(32'hb8e6dd13),
	.w7(32'h3b6be9c0),
	.w8(32'h3a97661d),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bee0208),
	.w1(32'h3c6889a8),
	.w2(32'h3bb89604),
	.w3(32'h3b4b800a),
	.w4(32'h3c24e472),
	.w5(32'h3c82ae44),
	.w6(32'h3afbfb21),
	.w7(32'hba6e7459),
	.w8(32'h3b8872b3),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3ca118),
	.w1(32'h3c79add2),
	.w2(32'h3b9cecd3),
	.w3(32'h3c0ec41e),
	.w4(32'h3c480942),
	.w5(32'h3c87a25b),
	.w6(32'h3c0dafbc),
	.w7(32'hbac4bea6),
	.w8(32'hbb003487),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba415c7),
	.w1(32'h3bbbd985),
	.w2(32'hbbea326b),
	.w3(32'h3c8f3a8f),
	.w4(32'h3b826f82),
	.w5(32'h3c17321d),
	.w6(32'h3b4a7d72),
	.w7(32'hbac9f923),
	.w8(32'hbb69cee1),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1709f6),
	.w1(32'h3c510524),
	.w2(32'hbb018c4a),
	.w3(32'h3ba93739),
	.w4(32'h3b91109f),
	.w5(32'h3c532303),
	.w6(32'h3a995df8),
	.w7(32'h3b3c1e2a),
	.w8(32'hbb8ed8a0),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9d07a0),
	.w1(32'h3bb176ce),
	.w2(32'h3c16b99a),
	.w3(32'h3b4ea042),
	.w4(32'hba3fb07e),
	.w5(32'hb9e56558),
	.w6(32'hb81ec2fa),
	.w7(32'h3af0fd11),
	.w8(32'h3bbcb107),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b017ec1),
	.w1(32'hb98f8d7d),
	.w2(32'h3c0c4cf0),
	.w3(32'h3bf81f44),
	.w4(32'hbb09f3ef),
	.w5(32'hbb775283),
	.w6(32'h3b44e56e),
	.w7(32'hbae83bed),
	.w8(32'hbb09a3d4),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab2f327),
	.w1(32'hbb364eed),
	.w2(32'hbb25425c),
	.w3(32'hbb2d8ccb),
	.w4(32'h394cccb2),
	.w5(32'hbb903914),
	.w6(32'h3a850476),
	.w7(32'h3b4aa903),
	.w8(32'h3b0152a2),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c96793d),
	.w1(32'h3c940bca),
	.w2(32'h3b872c4b),
	.w3(32'h3a4b6170),
	.w4(32'h3c2ab52f),
	.w5(32'h3c0a1b05),
	.w6(32'hbc0c1429),
	.w7(32'h3affcefe),
	.w8(32'h3c22d4cb),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c394754),
	.w1(32'h3bb55d51),
	.w2(32'hbaad8c54),
	.w3(32'hbaf65fe9),
	.w4(32'hbb2cf10b),
	.w5(32'hbbc29ab3),
	.w6(32'h3ace1e4f),
	.w7(32'h3b822610),
	.w8(32'hbab0e671),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa301a4),
	.w1(32'h3b923c16),
	.w2(32'h3bab7a90),
	.w3(32'hbc0fee59),
	.w4(32'h3adc21a2),
	.w5(32'hbb002a5f),
	.w6(32'hbb1558cb),
	.w7(32'h3b616866),
	.w8(32'h3b86b910),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1ea552),
	.w1(32'h3af2e70a),
	.w2(32'hbbeab3f6),
	.w3(32'hbb4b930d),
	.w4(32'hbc0ac192),
	.w5(32'hbc612382),
	.w6(32'h3a39c960),
	.w7(32'hbb1f73b1),
	.w8(32'hbbf701f6),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399fc557),
	.w1(32'h3bd0776a),
	.w2(32'h3b7b0e6e),
	.w3(32'hbbf32760),
	.w4(32'hba8f5037),
	.w5(32'h3b83b764),
	.w6(32'hbc2bb78f),
	.w7(32'h3a54d0dd),
	.w8(32'h3bc16eb5),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c3e1f5),
	.w1(32'h3c002a98),
	.w2(32'h3b11b5d8),
	.w3(32'h3b8e3f33),
	.w4(32'h3b7728a0),
	.w5(32'h3b328c56),
	.w6(32'h3bb0cf03),
	.w7(32'h3a4e43f2),
	.w8(32'hbad105eb),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1657c5),
	.w1(32'h3b062b21),
	.w2(32'h3bcd589f),
	.w3(32'h3ba7e389),
	.w4(32'hbaf9bdfa),
	.w5(32'hbb1d4c99),
	.w6(32'hba9baea5),
	.w7(32'hbc00ec15),
	.w8(32'h3b80e1f0),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b866eca),
	.w1(32'hbbd0e54e),
	.w2(32'hbb965be8),
	.w3(32'hbaecae51),
	.w4(32'h399c5c36),
	.w5(32'hbb480c2a),
	.w6(32'hbb940c59),
	.w7(32'h3a4c71dd),
	.w8(32'h398d84ef),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3f0a4f),
	.w1(32'hb9ccff7b),
	.w2(32'h3bb9243a),
	.w3(32'h3ad57eba),
	.w4(32'h3bb3e283),
	.w5(32'h3b33c376),
	.w6(32'h3bb3b9ad),
	.w7(32'h3c23d3f4),
	.w8(32'h3c0b8c81),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3169fc),
	.w1(32'h3a6ddc94),
	.w2(32'hb8b1df96),
	.w3(32'hbb0e2f7b),
	.w4(32'hbaa4ffb5),
	.w5(32'hbaa53c72),
	.w6(32'hb9d9519f),
	.w7(32'hbab4e87c),
	.w8(32'hbaa210b7),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c566a1e),
	.w1(32'h3c2b7066),
	.w2(32'h3bf53eb4),
	.w3(32'h3b850333),
	.w4(32'h3b05cce8),
	.w5(32'h3c9f7ce9),
	.w6(32'h3ae5fde7),
	.w7(32'h3a583482),
	.w8(32'h3c9116aa),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c61fe00),
	.w1(32'h3b013619),
	.w2(32'h3b0203fb),
	.w3(32'h3c03d60b),
	.w4(32'h3ba3f5f1),
	.w5(32'hbbe06994),
	.w6(32'h3c421491),
	.w7(32'hbaff5085),
	.w8(32'hbb38894b),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbef3323),
	.w1(32'hbc1bba08),
	.w2(32'h3b231c50),
	.w3(32'h3a342dd1),
	.w4(32'hbbc381a2),
	.w5(32'hba8615cb),
	.w6(32'h3acd424b),
	.w7(32'hbbacb360),
	.w8(32'hbbd93d6d),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b04f376),
	.w1(32'h3b1898fb),
	.w2(32'h3bf5b8ad),
	.w3(32'hbc1ab913),
	.w4(32'h3a94627e),
	.w5(32'h3cb70913),
	.w6(32'hbc164ff5),
	.w7(32'h3b06f399),
	.w8(32'h3c233b48),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9da22b),
	.w1(32'hbada20b4),
	.w2(32'h3bc1d34e),
	.w3(32'hbb09627e),
	.w4(32'hb9dcd0ff),
	.w5(32'hbac5b9f6),
	.w6(32'h3a3d4dc7),
	.w7(32'h3b4bab8d),
	.w8(32'hb99792ac),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4043aa),
	.w1(32'hbb4eec63),
	.w2(32'h3b657ff4),
	.w3(32'h3ba2d3ab),
	.w4(32'hbaf48cfa),
	.w5(32'h3b597e92),
	.w6(32'h3b3f9f7a),
	.w7(32'hbbb6b4f7),
	.w8(32'hbb7978bd),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a804bc7),
	.w1(32'hbbca5a0c),
	.w2(32'hba545e60),
	.w3(32'hbb983e89),
	.w4(32'h3b196df7),
	.w5(32'hbbf0e0b8),
	.w6(32'h3c023895),
	.w7(32'h3b540bb2),
	.w8(32'hbbb94ce9),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90ac436),
	.w1(32'h3bb1c741),
	.w2(32'h3c0bd9d0),
	.w3(32'hba904a6d),
	.w4(32'h3b970ad5),
	.w5(32'h3c052d5c),
	.w6(32'hbb89f471),
	.w7(32'hbb1040c3),
	.w8(32'hb9d3ea8d),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeff198),
	.w1(32'h3c1908b6),
	.w2(32'h3b866824),
	.w3(32'hbc3f479b),
	.w4(32'h3c9bee9d),
	.w5(32'h3a381201),
	.w6(32'hbad589ec),
	.w7(32'h3c5a3ade),
	.w8(32'h3b24f161),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7d5494),
	.w1(32'hbb360972),
	.w2(32'hbb3b5342),
	.w3(32'h3cb0b593),
	.w4(32'h3c009e02),
	.w5(32'hbc57cef9),
	.w6(32'hbad86b34),
	.w7(32'hbb7b82ad),
	.w8(32'hba944e52),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0871b1),
	.w1(32'h3b456f72),
	.w2(32'h3af1435b),
	.w3(32'h3c2d61d5),
	.w4(32'h3b694032),
	.w5(32'h3c40feaf),
	.w6(32'h3c01dc2b),
	.w7(32'hbb91869f),
	.w8(32'h3c22927a),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baea338),
	.w1(32'h3c849273),
	.w2(32'h3c4e3a2f),
	.w3(32'hbb762d33),
	.w4(32'h3c95e206),
	.w5(32'h3c51de10),
	.w6(32'h3b2968da),
	.w7(32'h3bf4f6f5),
	.w8(32'h3bd48280),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd2af14),
	.w1(32'hbc09f892),
	.w2(32'hbb84e031),
	.w3(32'h3bc8659b),
	.w4(32'hbbe99cbd),
	.w5(32'hbbd2730a),
	.w6(32'h3bce4eaf),
	.w7(32'hbc0066d4),
	.w8(32'hbb90830a),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabd47d8),
	.w1(32'hbb57ccf6),
	.w2(32'h38f32b85),
	.w3(32'h39f9f70f),
	.w4(32'h3b7f0438),
	.w5(32'h3be41284),
	.w6(32'hb9e16559),
	.w7(32'h3ad6b333),
	.w8(32'hb99ad435),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a88bc99),
	.w1(32'h3b104c1d),
	.w2(32'h3c070b4d),
	.w3(32'hba0b9a4d),
	.w4(32'h3a9a35a4),
	.w5(32'h3b9da263),
	.w6(32'hbb29a314),
	.w7(32'hbb65907a),
	.w8(32'h3b147b80),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba5f0a3),
	.w1(32'h3ae0b7d7),
	.w2(32'h3b8a25c4),
	.w3(32'h3b3c4894),
	.w4(32'hbb4a5054),
	.w5(32'h3b2d13d5),
	.w6(32'hbbaff117),
	.w7(32'hbc4284d1),
	.w8(32'hbb49ffa9),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4b2a66),
	.w1(32'hbba59fe7),
	.w2(32'hba60deeb),
	.w3(32'hb85a955b),
	.w4(32'h3a839585),
	.w5(32'hbbe8dda3),
	.w6(32'hbb787fde),
	.w7(32'hbbd0b0d7),
	.w8(32'hbb3d2bf4),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbd46ec),
	.w1(32'hbb04971e),
	.w2(32'hbc22dfc9),
	.w3(32'hbabf1513),
	.w4(32'hbc4eb172),
	.w5(32'h3ab44da0),
	.w6(32'hbc8066b7),
	.w7(32'hbc6a465f),
	.w8(32'hbb41d20b),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc60c067),
	.w1(32'hbbbb8d2d),
	.w2(32'hbb1b0648),
	.w3(32'hbca2306f),
	.w4(32'hbc1c74c5),
	.w5(32'hbc41c5a2),
	.w6(32'hbba87a04),
	.w7(32'hbbb964f1),
	.w8(32'hbc10cf81),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc23f6f3),
	.w1(32'hba3d6b32),
	.w2(32'h3b20e732),
	.w3(32'hbc93344c),
	.w4(32'hbaff97f5),
	.w5(32'hbbc1cc5d),
	.w6(32'hbc515b45),
	.w7(32'hbb4c2f09),
	.w8(32'hbb5ccf3e),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7c0c83),
	.w1(32'h3b458b4a),
	.w2(32'h3c3ace64),
	.w3(32'hbb6d70e1),
	.w4(32'hbbc4dfbe),
	.w5(32'h3a2e34f6),
	.w6(32'hba1d725c),
	.w7(32'h3b4bbba7),
	.w8(32'hb78c9ea2),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8e9510),
	.w1(32'h3c731cd8),
	.w2(32'h3bda7f13),
	.w3(32'h3c8002f5),
	.w4(32'h3ab966de),
	.w5(32'h3c3f8cd3),
	.w6(32'hba9d7210),
	.w7(32'hbab1ae47),
	.w8(32'h3c3005eb),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7f911d),
	.w1(32'h3be3ba49),
	.w2(32'h3c1f32ed),
	.w3(32'h39234c39),
	.w4(32'hbbb824be),
	.w5(32'hbbf34652),
	.w6(32'hbb6eb1c3),
	.w7(32'hbc061edb),
	.w8(32'hbb2cc087),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa685e6),
	.w1(32'h3b1bf2e8),
	.w2(32'hba8181df),
	.w3(32'hbb6a09eb),
	.w4(32'h3ba38597),
	.w5(32'hbb5f6b70),
	.w6(32'hbbd15505),
	.w7(32'hbb6a3f04),
	.w8(32'h3a97e5a3),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b65de0e),
	.w1(32'h3ba0be3a),
	.w2(32'h3b4883c7),
	.w3(32'h3c414b6f),
	.w4(32'h3b0fbd4a),
	.w5(32'h3b04cb2d),
	.w6(32'h3c6d2665),
	.w7(32'h3bd16986),
	.w8(32'h3b20379d),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb688b30),
	.w1(32'hba7ba372),
	.w2(32'h3b496a3d),
	.w3(32'h39b49fdf),
	.w4(32'h3c129aa7),
	.w5(32'h3a89f3da),
	.w6(32'hba12cc22),
	.w7(32'hb9cb1c5d),
	.w8(32'h3c01c778),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb32e225),
	.w1(32'h3bb85b8a),
	.w2(32'h3c1a3ed9),
	.w3(32'hbc088c82),
	.w4(32'hbbd66be5),
	.w5(32'h3bf05ad6),
	.w6(32'hb8256c44),
	.w7(32'h3b796e79),
	.w8(32'h3bc13f2a),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8e4d78),
	.w1(32'hbbb16df7),
	.w2(32'h3bb083b0),
	.w3(32'h3c8a82f8),
	.w4(32'hbabb4d53),
	.w5(32'hbaf50296),
	.w6(32'h3bad482c),
	.w7(32'hbc004eb4),
	.w8(32'hbb406fa9),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc11038),
	.w1(32'h3b3fe57b),
	.w2(32'h3ac63dcd),
	.w3(32'hbbedbd44),
	.w4(32'h3bb20fac),
	.w5(32'h3b9c6d96),
	.w6(32'hbc17c111),
	.w7(32'h3bbad685),
	.w8(32'hbacc8c4c),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9e6101),
	.w1(32'h3b90966f),
	.w2(32'h3b694315),
	.w3(32'hb9d69f84),
	.w4(32'h3ae98b57),
	.w5(32'h3c3c3c39),
	.w6(32'hb92bf425),
	.w7(32'h3a746269),
	.w8(32'h3c08b931),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7202ff),
	.w1(32'h3b274509),
	.w2(32'hbb688cfd),
	.w3(32'h3a3214d7),
	.w4(32'hbc223a6d),
	.w5(32'hbc2d1d9e),
	.w6(32'hbaffe140),
	.w7(32'hbc0b83f2),
	.w8(32'hbb1aac36),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2aa42a),
	.w1(32'h3a881272),
	.w2(32'h3b52a860),
	.w3(32'hba9c74a7),
	.w4(32'h3afb083c),
	.w5(32'h3a61d5b5),
	.w6(32'hbb79a011),
	.w7(32'hbbb16b4a),
	.w8(32'h3b4e6d31),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a83edb3),
	.w1(32'hbaefc318),
	.w2(32'hbae3826d),
	.w3(32'h3a4119a8),
	.w4(32'hbbadafc7),
	.w5(32'h3bc9b60a),
	.w6(32'h3bbee7c4),
	.w7(32'hbbb2b507),
	.w8(32'h3b9f8a9e),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc730ebe),
	.w1(32'h3c7d9851),
	.w2(32'h3c84b919),
	.w3(32'hbc962055),
	.w4(32'h3b928427),
	.w5(32'h3c55f71f),
	.w6(32'hbc9fc4ef),
	.w7(32'h3b8f398d),
	.w8(32'h3c292d63),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c439683),
	.w1(32'h3aa7d986),
	.w2(32'hbb8a53c6),
	.w3(32'h3b9bebef),
	.w4(32'h3b59758d),
	.w5(32'hbbe984aa),
	.w6(32'hbbbeacdf),
	.w7(32'h3b273616),
	.w8(32'h3a177322),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be37dab),
	.w1(32'h3bca70ac),
	.w2(32'h3bae3732),
	.w3(32'h3bf8dd69),
	.w4(32'h3caba237),
	.w5(32'hb9d83366),
	.w6(32'hbb8689dd),
	.w7(32'h3bacb81d),
	.w8(32'hbba3be4f),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8c6e9d),
	.w1(32'h3aa3bd18),
	.w2(32'h3a1cd89c),
	.w3(32'h3b75f84f),
	.w4(32'hb9f0e466),
	.w5(32'hb9333183),
	.w6(32'h3bb0e5ff),
	.w7(32'hbb9f4501),
	.w8(32'h39f0c019),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1411a8),
	.w1(32'h3baaa66b),
	.w2(32'hba6c5385),
	.w3(32'hb8e141ee),
	.w4(32'h3c428d9f),
	.w5(32'hbb356e5d),
	.w6(32'hbaddcef5),
	.w7(32'h3b99f796),
	.w8(32'hbb12ff0d),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b36d22b),
	.w1(32'h3a0d57e8),
	.w2(32'h3ad03667),
	.w3(32'h3b5bbf19),
	.w4(32'h39647377),
	.w5(32'hbb16238d),
	.w6(32'h3a005253),
	.w7(32'h3b0f5052),
	.w8(32'hbb00fc53),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b493f8f),
	.w1(32'hbb04b990),
	.w2(32'h3b35e9e4),
	.w3(32'h3c657780),
	.w4(32'h3b42237b),
	.w5(32'h3b092e96),
	.w6(32'h3bd483a0),
	.w7(32'h3c076069),
	.w8(32'h3b6152b6),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba339c4f),
	.w1(32'h3c5f3040),
	.w2(32'h3c988f53),
	.w3(32'hbb6449df),
	.w4(32'h3c28415e),
	.w5(32'h3cc079a6),
	.w6(32'hbb83bdac),
	.w7(32'hba61da49),
	.w8(32'h3c688297),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c205b1b),
	.w1(32'hbbe2b7d0),
	.w2(32'hbc54566f),
	.w3(32'h3c3837e6),
	.w4(32'hbbda799a),
	.w5(32'h3b6c6758),
	.w6(32'h3ca178a4),
	.w7(32'h3b8dd1ad),
	.w8(32'h39837b3e),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3708c1),
	.w1(32'h3b5c2aa0),
	.w2(32'h392c07f0),
	.w3(32'h3c22834c),
	.w4(32'hb881f6c5),
	.w5(32'hbabb6d83),
	.w6(32'hbc229c0f),
	.w7(32'hbbb2a2a3),
	.w8(32'h3a4302e5),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdcdf21),
	.w1(32'h3c24db06),
	.w2(32'h3c19a4aa),
	.w3(32'h3a082b07),
	.w4(32'h3af58c52),
	.w5(32'hbb88c5b1),
	.w6(32'hbbb60f76),
	.w7(32'h3a8c7e74),
	.w8(32'hba69b8e3),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c949c8a),
	.w1(32'h3c26b261),
	.w2(32'h3b870493),
	.w3(32'h3c19662a),
	.w4(32'h3bec6993),
	.w5(32'h3b416bd5),
	.w6(32'h3b11a42a),
	.w7(32'h3b369fa2),
	.w8(32'h3b9f6b8c),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b905e47),
	.w1(32'hbace49b4),
	.w2(32'hbaf59803),
	.w3(32'h3bd5d9ee),
	.w4(32'h3be0b3dc),
	.w5(32'hbaf086c1),
	.w6(32'h3ad7f4b7),
	.w7(32'h3a90381b),
	.w8(32'hbaa15e69),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h379136b7),
	.w1(32'h3b86448b),
	.w2(32'hbacd5935),
	.w3(32'hbb8bbf34),
	.w4(32'h3a896620),
	.w5(32'hbbd59c4a),
	.w6(32'h3b3653ba),
	.w7(32'hbb51f581),
	.w8(32'hba28c9c1),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f2080f),
	.w1(32'h3c10745e),
	.w2(32'h3c0da55f),
	.w3(32'h3bea1a19),
	.w4(32'h3b74aa71),
	.w5(32'h3c3910f0),
	.w6(32'h3b8d1b65),
	.w7(32'h3a815496),
	.w8(32'h3c35805d),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beb6262),
	.w1(32'hbb840e28),
	.w2(32'hbabfbdfd),
	.w3(32'hbb9f6aa5),
	.w4(32'hbb266c9a),
	.w5(32'hba8d825e),
	.w6(32'h3b86a7f3),
	.w7(32'h3b3fff30),
	.w8(32'hbaf58a27),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3b353e),
	.w1(32'h3b8e99c1),
	.w2(32'h3ba03790),
	.w3(32'hbbad195f),
	.w4(32'h3b5b2bfa),
	.w5(32'h3ae30bc0),
	.w6(32'hb7b6ee3c),
	.w7(32'h3c12df02),
	.w8(32'hba60520b),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c059812),
	.w1(32'h3b56e8bf),
	.w2(32'h3c2c1033),
	.w3(32'h3be50d2b),
	.w4(32'hb9f318e9),
	.w5(32'h3cf37241),
	.w6(32'hbb56f97f),
	.w7(32'hbb4e558c),
	.w8(32'h3c6e67b7),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd03d0c),
	.w1(32'h3b447eb2),
	.w2(32'hbb14e99e),
	.w3(32'hbc1f87f6),
	.w4(32'h3ae77142),
	.w5(32'hbba205b3),
	.w6(32'hbbc41522),
	.w7(32'hbbaeddfd),
	.w8(32'hbaa27d1a),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8412e5),
	.w1(32'h3bf6a155),
	.w2(32'hbb95c8a8),
	.w3(32'h39e4dc82),
	.w4(32'h3b30c7e5),
	.w5(32'h3b7db668),
	.w6(32'h3ba0032d),
	.w7(32'h3bfdb955),
	.w8(32'h3c17e197),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2e3aec),
	.w1(32'hbc2a3cf3),
	.w2(32'hbb5098b8),
	.w3(32'h3c4219fc),
	.w4(32'hbba7ffff),
	.w5(32'hbc720604),
	.w6(32'h3bd38d6c),
	.w7(32'hbc08392c),
	.w8(32'hbc1f0b44),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1bf462),
	.w1(32'hbbd54667),
	.w2(32'hbb9f0edf),
	.w3(32'hbcaa2226),
	.w4(32'hbb8d897d),
	.w5(32'hbc0c07d2),
	.w6(32'hbc7f6c34),
	.w7(32'hbc246a10),
	.w8(32'hbbdb4d94),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9ca09f),
	.w1(32'hbbea9f99),
	.w2(32'h3a10a4cc),
	.w3(32'hbb0120e1),
	.w4(32'hbbc7920c),
	.w5(32'hbc06d8e2),
	.w6(32'hbbd6a06a),
	.w7(32'hbbb73630),
	.w8(32'hb816c638),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0ad2a1),
	.w1(32'h3c8dad6c),
	.w2(32'h3c09eebc),
	.w3(32'hbc875928),
	.w4(32'h3c5ba874),
	.w5(32'hbbab5acb),
	.w6(32'hbc7a6670),
	.w7(32'hba2603b6),
	.w8(32'hb8ab6530),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3badb00e),
	.w1(32'h3b1069b1),
	.w2(32'h3bc1e1be),
	.w3(32'h3c0d8efd),
	.w4(32'h3ab0e469),
	.w5(32'h3c045c2d),
	.w6(32'h3c555c4c),
	.w7(32'hbb3aacd0),
	.w8(32'h3bcf073f),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbb14df),
	.w1(32'hbb87a64e),
	.w2(32'h3c32a41f),
	.w3(32'h3c5505b4),
	.w4(32'hbbafa49f),
	.w5(32'h3b4b1176),
	.w6(32'h3c1158a5),
	.w7(32'hbbd18351),
	.w8(32'hbc2056a5),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule