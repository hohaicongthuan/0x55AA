module layer_8_featuremap_119(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4a23d0),
	.w1(32'hbaf17eb1),
	.w2(32'h3bb88dbc),
	.w3(32'h3adf8392),
	.w4(32'hbb9319ef),
	.w5(32'hbb8a97a5),
	.w6(32'h36b45c58),
	.w7(32'hbb863fcd),
	.w8(32'hbc4158b8),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf6b3f1),
	.w1(32'h3bfadd6e),
	.w2(32'hba9f5586),
	.w3(32'h3c4ddffe),
	.w4(32'hbc1b5065),
	.w5(32'hbc5485a1),
	.w6(32'hbb19ec33),
	.w7(32'hbc1ac974),
	.w8(32'h3a8b009c),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1e6047),
	.w1(32'hba575d43),
	.w2(32'h3c057b2c),
	.w3(32'hbb3d46e3),
	.w4(32'h3bd762f9),
	.w5(32'hbc36b42d),
	.w6(32'h3b5d10ed),
	.w7(32'h3cb94cfa),
	.w8(32'hbc7bb103),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc59eab),
	.w1(32'hbbc671b8),
	.w2(32'hbc525425),
	.w3(32'hb80abdbd),
	.w4(32'hbb61ed00),
	.w5(32'h3b8258dd),
	.w6(32'h3aa74ce8),
	.w7(32'hbc56ef4a),
	.w8(32'hbbe3a2dd),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5e3936),
	.w1(32'h3aaed9e8),
	.w2(32'h3c19cf51),
	.w3(32'hbb912d23),
	.w4(32'hbc05355a),
	.w5(32'hbc149671),
	.w6(32'h3c77deb8),
	.w7(32'h3bd2b539),
	.w8(32'hbcad6038),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb319271),
	.w1(32'hbc6e0412),
	.w2(32'h3c2ad65e),
	.w3(32'hbc272e66),
	.w4(32'hbb4e7182),
	.w5(32'h3bfd3f86),
	.w6(32'hbbed940d),
	.w7(32'h3bafa8b0),
	.w8(32'h3bd7602c),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc387c1a),
	.w1(32'h3bfadea4),
	.w2(32'h3b8bef7b),
	.w3(32'hbb51a4e3),
	.w4(32'hba9e7cfe),
	.w5(32'h3b6ac477),
	.w6(32'h3c09784e),
	.w7(32'hbb5a7946),
	.w8(32'hbc8c2621),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc046785),
	.w1(32'h3c32abcc),
	.w2(32'h3cc27e8a),
	.w3(32'h3cab9a76),
	.w4(32'hbb440241),
	.w5(32'hbb54e3c3),
	.w6(32'h3c3877dc),
	.w7(32'h3c2360a2),
	.w8(32'hbc844f25),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcba7657),
	.w1(32'h3bf34e12),
	.w2(32'h3c814ac1),
	.w3(32'hbb7984d9),
	.w4(32'h3ca3a137),
	.w5(32'h3b595e74),
	.w6(32'h3bcdbac5),
	.w7(32'h3be9240b),
	.w8(32'hb9defca1),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc465f90),
	.w1(32'hbbda6d8a),
	.w2(32'hbbae2bfb),
	.w3(32'hbb4dedeb),
	.w4(32'h3acc863e),
	.w5(32'hbb2322b2),
	.w6(32'hbbd9ba55),
	.w7(32'h3c07a5f1),
	.w8(32'h3d1434a2),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0a798b),
	.w1(32'h3ca7eeb5),
	.w2(32'h3cb54d83),
	.w3(32'hbc72d5ab),
	.w4(32'h3c8d8166),
	.w5(32'hbc1af780),
	.w6(32'hbc52f632),
	.w7(32'h3d62f721),
	.w8(32'hbd13ab11),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb0dca3),
	.w1(32'hb8bd7cbe),
	.w2(32'h3c10119b),
	.w3(32'hbb168c2c),
	.w4(32'hbc47f6bc),
	.w5(32'hbc8bff18),
	.w6(32'h3cce057a),
	.w7(32'hbc1c3bdc),
	.w8(32'hbd05785d),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc83c7b7),
	.w1(32'hba2b63e1),
	.w2(32'h394bfde0),
	.w3(32'h39c96b42),
	.w4(32'h3955a29a),
	.w5(32'hb91d6cab),
	.w6(32'hbb80d2ec),
	.w7(32'h3b1ad9a4),
	.w8(32'h3b226cfe),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a73fec),
	.w1(32'h398f4163),
	.w2(32'h3a47c2f3),
	.w3(32'h398c2a14),
	.w4(32'h3a3c8fdb),
	.w5(32'h3a5f6e11),
	.w6(32'h3a08951a),
	.w7(32'h39b8e22f),
	.w8(32'h395f5ca4),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37882a77),
	.w1(32'h389b0923),
	.w2(32'h391c8c5e),
	.w3(32'h3890071f),
	.w4(32'h39016347),
	.w5(32'h3922ecaf),
	.w6(32'h38c1709d),
	.w7(32'h39411291),
	.w8(32'h39407c90),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6d6dd4),
	.w1(32'h3a6fc40e),
	.w2(32'h3a72bc6b),
	.w3(32'h3a9a747f),
	.w4(32'h3a8944b1),
	.w5(32'h3a3e3f8b),
	.w6(32'h3a7d4e1e),
	.w7(32'h3a807b32),
	.w8(32'h3a63bec5),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba44b14d),
	.w1(32'hba5be86d),
	.w2(32'hb9f0f5b9),
	.w3(32'h3a54d4fa),
	.w4(32'hb8cba435),
	.w5(32'hb9073d62),
	.w6(32'h3a8a4ad7),
	.w7(32'h3a4ae89e),
	.w8(32'h3a144ef1),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b21bf6b),
	.w1(32'h3aaa6437),
	.w2(32'h3b6426af),
	.w3(32'h3b886293),
	.w4(32'h3b15affe),
	.w5(32'h3b5a99bc),
	.w6(32'h3b6bc3ec),
	.w7(32'h3b06ec4f),
	.w8(32'h3b0fcf40),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c58fef4),
	.w1(32'h3c4e7c56),
	.w2(32'h3c08987a),
	.w3(32'h3c3c9f06),
	.w4(32'h3c032b81),
	.w5(32'h3a76b098),
	.w6(32'h3bea8107),
	.w7(32'h39169478),
	.w8(32'hbba885b4),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c04a2d8),
	.w1(32'h3be78e3f),
	.w2(32'h3bd243d7),
	.w3(32'h3c1a9af5),
	.w4(32'h3c17ecd8),
	.w5(32'h3bba61b7),
	.w6(32'hba00ee65),
	.w7(32'hba0b17d6),
	.w8(32'hbb5d30f1),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb82905a5),
	.w1(32'h3a0b49ca),
	.w2(32'h3b336585),
	.w3(32'hbb299624),
	.w4(32'hbae77725),
	.w5(32'h3ac7872f),
	.w6(32'hbaa682b4),
	.w7(32'hbb04838b),
	.w8(32'hba8251d0),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2662bf),
	.w1(32'h383cdd99),
	.w2(32'h3b71151e),
	.w3(32'h3b2a84ab),
	.w4(32'h3a36a0a2),
	.w5(32'h3ba65cf5),
	.w6(32'h3b2573a4),
	.w7(32'h3b040e1f),
	.w8(32'h3b862915),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2343c5),
	.w1(32'h3bb90791),
	.w2(32'h3ad92f04),
	.w3(32'h3b84a1a5),
	.w4(32'h3bf99895),
	.w5(32'hbaa168ef),
	.w6(32'hbbda58c2),
	.w7(32'hbc042692),
	.w8(32'hbc432a07),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac7883c),
	.w1(32'hbadf16bd),
	.w2(32'h39e252eb),
	.w3(32'hb90f53c7),
	.w4(32'h3ae20c48),
	.w5(32'h3b106a30),
	.w6(32'h3a919df2),
	.w7(32'h3aeecbaa),
	.w8(32'h3b11a441),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b12fccd),
	.w1(32'h3a87a073),
	.w2(32'h3ab7183c),
	.w3(32'h3ab073f1),
	.w4(32'h39957b46),
	.w5(32'h399e4c47),
	.w6(32'h3b112341),
	.w7(32'h3abbbef7),
	.w8(32'h3ac25dad),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e9fd31),
	.w1(32'h3b1d7ac4),
	.w2(32'h3b5cf811),
	.w3(32'h3afd8988),
	.w4(32'h3b99ed10),
	.w5(32'h3ac95a85),
	.w6(32'hbb80b8e5),
	.w7(32'hbb37de5f),
	.w8(32'hbb51650f),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba757762),
	.w1(32'hba68ac15),
	.w2(32'hba6840d1),
	.w3(32'hba85a6ab),
	.w4(32'hbaa0e1a8),
	.w5(32'hba538a9d),
	.w6(32'hbae1e692),
	.w7(32'hbae0b306),
	.w8(32'hba16cfaa),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc166d1),
	.w1(32'h3bcc33ce),
	.w2(32'h3c09afca),
	.w3(32'h3ce64b30),
	.w4(32'h3befe1e2),
	.w5(32'h3c9f3bc5),
	.w6(32'h3c87ea96),
	.w7(32'hbcce92f4),
	.w8(32'hbcc0f074),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b396709),
	.w1(32'h3b22cfad),
	.w2(32'h3b059704),
	.w3(32'h3b25c7eb),
	.w4(32'h3ada322e),
	.w5(32'h3a1d0c64),
	.w6(32'h39b8d142),
	.w7(32'hba5f4487),
	.w8(32'hbaa97a7e),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af13af4),
	.w1(32'h3ac7cbe7),
	.w2(32'h3b4c33d6),
	.w3(32'h3b02cd27),
	.w4(32'h3ae5b3ae),
	.w5(32'h3b253e11),
	.w6(32'h3b0d6fb6),
	.w7(32'h3acda15d),
	.w8(32'h3b0952dd),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9eeae3),
	.w1(32'hbb9f2713),
	.w2(32'hbb13d947),
	.w3(32'hbb9b0e39),
	.w4(32'hbbcc35d3),
	.w5(32'hbb2ea39b),
	.w6(32'hbb469d8b),
	.w7(32'hbb68f3d6),
	.w8(32'hb94a919e),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9d01fd),
	.w1(32'h3a9c41e8),
	.w2(32'h3b0cf5ed),
	.w3(32'h3ac89ac8),
	.w4(32'h3a3ef127),
	.w5(32'h3a1e74e2),
	.w6(32'hb90596ed),
	.w7(32'hba6b8cd0),
	.w8(32'hb98730f8),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97f2e85),
	.w1(32'hb9018e0e),
	.w2(32'hb8bfa109),
	.w3(32'hb9565d7a),
	.w4(32'hb178fb40),
	.w5(32'hb82ed0ff),
	.w6(32'hb7f714c3),
	.w7(32'h393cc8a5),
	.w8(32'h38e927eb),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8dede9c),
	.w1(32'hb8301965),
	.w2(32'hb8beea38),
	.w3(32'hb85c8a44),
	.w4(32'h383f2128),
	.w5(32'hb789abbd),
	.w6(32'hb8abace9),
	.w7(32'h378a7e4d),
	.w8(32'hb7fa95bb),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae9740f),
	.w1(32'hbb61f1c3),
	.w2(32'hbada776f),
	.w3(32'hba0bd9d8),
	.w4(32'hbaa1cda9),
	.w5(32'h39bf21f7),
	.w6(32'hba389b32),
	.w7(32'hbad0d53c),
	.w8(32'hb958f73d),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a946a40),
	.w1(32'h3b728618),
	.w2(32'h3b206480),
	.w3(32'h3aa9ed13),
	.w4(32'h3aec5584),
	.w5(32'h3a2dc153),
	.w6(32'h38c4ec3f),
	.w7(32'h39c49084),
	.w8(32'hba06dcae),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389b2351),
	.w1(32'h398564f8),
	.w2(32'h391b0d34),
	.w3(32'h3a1a9ed7),
	.w4(32'h3a10a50c),
	.w5(32'h3999d71c),
	.w6(32'h39b13792),
	.w7(32'h3992873f),
	.w8(32'h39a2c179),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afa5c93),
	.w1(32'h3b5240c7),
	.w2(32'h3b8b6bb5),
	.w3(32'h3a861807),
	.w4(32'h3b0f1f4f),
	.w5(32'h3b2b6c56),
	.w6(32'hb9e37430),
	.w7(32'hba45aca2),
	.w8(32'h3a028699),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38535b74),
	.w1(32'h39e630e1),
	.w2(32'hb9a4b05d),
	.w3(32'h3987dab5),
	.w4(32'h3a19caaf),
	.w5(32'h39cff354),
	.w6(32'h38a13439),
	.w7(32'h39d1efe4),
	.w8(32'h37c30f74),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89ebd79),
	.w1(32'hb9485b33),
	.w2(32'hb9ec74fe),
	.w3(32'h39282b13),
	.w4(32'h3804833e),
	.w5(32'hb8b5a699),
	.w6(32'hb706ecaf),
	.w7(32'hb8c02b20),
	.w8(32'hb98be210),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb919d6),
	.w1(32'h3b5dfa85),
	.w2(32'h3bd552fd),
	.w3(32'h3babd96b),
	.w4(32'h3b155354),
	.w5(32'h3b9c8b1d),
	.w6(32'h3ab5253e),
	.w7(32'hba1226f5),
	.w8(32'h3b7e69d5),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e7d8c8),
	.w1(32'h39c35294),
	.w2(32'hba1686c9),
	.w3(32'h3a708e89),
	.w4(32'h39e22ae1),
	.w5(32'hba1f2f55),
	.w6(32'h39dce173),
	.w7(32'hba6e72b4),
	.w8(32'hbabb0bd1),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b53208),
	.w1(32'hb8fd9d69),
	.w2(32'hb98b9d49),
	.w3(32'hb67754e9),
	.w4(32'hb836697f),
	.w5(32'hb9039907),
	.w6(32'h38c9877f),
	.w7(32'h38336840),
	.w8(32'hb89979fc),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8a7d72),
	.w1(32'h3a595d96),
	.w2(32'h3a246a6d),
	.w3(32'h3af5772a),
	.w4(32'h3a69034c),
	.w5(32'h39a86556),
	.w6(32'h3899bdcf),
	.w7(32'hba768a11),
	.w8(32'hba59083e),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b23bb3f),
	.w1(32'h3b18becb),
	.w2(32'h3b3d4d83),
	.w3(32'h3b76522b),
	.w4(32'h3afb501c),
	.w5(32'h3ab4a612),
	.w6(32'h38728071),
	.w7(32'hbb2b800e),
	.w8(32'hbb464f3a),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388c296b),
	.w1(32'hbaa38ccd),
	.w2(32'hbabbeebf),
	.w3(32'hba88ba4b),
	.w4(32'hbadbaf7b),
	.w5(32'hbb088d36),
	.w6(32'hba02fd59),
	.w7(32'hbaa62569),
	.w8(32'hbab49825),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb848bab6),
	.w1(32'hb79450e2),
	.w2(32'hb83ffb46),
	.w3(32'hb785f7f3),
	.w4(32'h37a78c47),
	.w5(32'hb7d10b12),
	.w6(32'hb785929f),
	.w7(32'h37979b2d),
	.w8(32'hb79aeed9),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8d33d1),
	.w1(32'h3beb799c),
	.w2(32'h3b907436),
	.w3(32'h3be5683a),
	.w4(32'h3c026e91),
	.w5(32'h3b351ec0),
	.w6(32'h3b5ac375),
	.w7(32'h3aa00467),
	.w8(32'hbb8ddd39),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b277f79),
	.w1(32'h3aa3319e),
	.w2(32'h3aa4a1bc),
	.w3(32'h3b2a063d),
	.w4(32'h3ab67935),
	.w5(32'h3aa93636),
	.w6(32'h3b15a2b8),
	.w7(32'h3a8cd532),
	.w8(32'h3aa802b9),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b639eb3),
	.w1(32'h3b2ee7f0),
	.w2(32'h3b0667c4),
	.w3(32'h3b7711ad),
	.w4(32'h3b366e7e),
	.w5(32'h3ace0e64),
	.w6(32'h3ac011c2),
	.w7(32'h393228db),
	.w8(32'h388b2c3e),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a858adc),
	.w1(32'hba844ae0),
	.w2(32'h3b4bb8ef),
	.w3(32'h39828031),
	.w4(32'hbb22445f),
	.w5(32'h3a3e8307),
	.w6(32'hbb06c9d9),
	.w7(32'hbb93f3c9),
	.w8(32'hba3f0e58),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3c753e),
	.w1(32'h3c4a978e),
	.w2(32'h3c1f94e0),
	.w3(32'h3c9bada6),
	.w4(32'h3c900c55),
	.w5(32'h3c422e56),
	.w6(32'h3b88908b),
	.w7(32'hb939cac6),
	.w8(32'hbbc06553),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0f1ef4),
	.w1(32'h3a6ef0b5),
	.w2(32'hbb30fd52),
	.w3(32'h3bdaf3f2),
	.w4(32'h3baa62da),
	.w5(32'hb93f4514),
	.w6(32'h3a805535),
	.w7(32'h39631ad0),
	.w8(32'hbb94ae41),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af68798),
	.w1(32'h3aa13ffb),
	.w2(32'h3a99f22a),
	.w3(32'h3b344ba9),
	.w4(32'h3acf8bb4),
	.w5(32'h3a9c830e),
	.w6(32'h3b7b9f29),
	.w7(32'h3afdc7ff),
	.w8(32'h3ad85aa2),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d320e5),
	.w1(32'h381a9ad7),
	.w2(32'hb7d922a6),
	.w3(32'hb84e0fa4),
	.w4(32'h38c04789),
	.w5(32'h38423df7),
	.w6(32'hb7f6717f),
	.w7(32'h38da9f1b),
	.w8(32'h38b4c3db),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4629d0),
	.w1(32'h3b92fe83),
	.w2(32'h3ba86395),
	.w3(32'h3ba69ed6),
	.w4(32'h3b83e6d1),
	.w5(32'h3b107583),
	.w6(32'h3a8c72db),
	.w7(32'hbae36e58),
	.w8(32'hb9a315d6),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94ef3b5),
	.w1(32'hbaea9444),
	.w2(32'hba3c2035),
	.w3(32'h3b2485d3),
	.w4(32'h3a22d04c),
	.w5(32'h3a502cb7),
	.w6(32'h3a7e70d0),
	.w7(32'hba6b7ec5),
	.w8(32'hb97c1a34),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeb0cb2),
	.w1(32'h3a97956b),
	.w2(32'h3af9b735),
	.w3(32'h3b95a684),
	.w4(32'h3b665756),
	.w5(32'h3b6535a2),
	.w6(32'h3ab77852),
	.w7(32'h3a9f2094),
	.w8(32'h3b2983fe),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af6850f),
	.w1(32'h3b1636cc),
	.w2(32'h3b045edf),
	.w3(32'h3b5c1193),
	.w4(32'h3b46dba0),
	.w5(32'h3b076b2c),
	.w6(32'h3a79ddd5),
	.w7(32'hba5e77ef),
	.w8(32'hbb080f5d),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8652bb),
	.w1(32'h3a9de004),
	.w2(32'h3a727d00),
	.w3(32'h3b125dea),
	.w4(32'h3b1f8148),
	.w5(32'h3aacb2cc),
	.w6(32'h3afacffd),
	.w7(32'h3aabf1dc),
	.w8(32'h39582a96),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a12f8d8),
	.w1(32'h39b0ce39),
	.w2(32'h362b3736),
	.w3(32'h3a94b718),
	.w4(32'h3a5a566e),
	.w5(32'h39dafcf8),
	.w6(32'h3aa9a6c3),
	.w7(32'h3a8b099c),
	.w8(32'h3a51f984),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3971c56e),
	.w1(32'h393a952e),
	.w2(32'h3981501b),
	.w3(32'h3a14a829),
	.w4(32'h3a1a80e8),
	.w5(32'h39ddec84),
	.w6(32'h39d5c724),
	.w7(32'h3987a4a3),
	.w8(32'h38ea7c59),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9799b7),
	.w1(32'h3b645773),
	.w2(32'h3b828aa0),
	.w3(32'h3b8f9ba3),
	.w4(32'h3b1a4ece),
	.w5(32'h3b0dea69),
	.w6(32'h3ac637e9),
	.w7(32'hb9fb2921),
	.w8(32'h3a3a95dc),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a08cb36),
	.w1(32'h39fab525),
	.w2(32'hb7bc4c42),
	.w3(32'h3b140c25),
	.w4(32'h3ae9b05d),
	.w5(32'h3ac962c1),
	.w6(32'h3b10b750),
	.w7(32'h3b0b2c18),
	.w8(32'h39f237a1),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8a6e0e),
	.w1(32'hba11ea75),
	.w2(32'hba64d214),
	.w3(32'hb9f8c208),
	.w4(32'h390c841b),
	.w5(32'hba1d82ee),
	.w6(32'hba42f182),
	.w7(32'h38908975),
	.w8(32'hba476773),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba92aebe),
	.w1(32'hb9d8abb5),
	.w2(32'hb943bba3),
	.w3(32'h3a245449),
	.w4(32'h3ac5b878),
	.w5(32'h3a9a93fa),
	.w6(32'hb79702a0),
	.w7(32'h39b39cb7),
	.w8(32'h39726536),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3f4b05),
	.w1(32'h3b00f4a0),
	.w2(32'h3b61ce1d),
	.w3(32'h3b622519),
	.w4(32'h3b429ba8),
	.w5(32'h3b63097b),
	.w6(32'h3b0be6f9),
	.w7(32'h3ac855be),
	.w8(32'h3abfd648),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb974b929),
	.w1(32'hbab116ed),
	.w2(32'hba5f8575),
	.w3(32'hba0914e7),
	.w4(32'hbabaea44),
	.w5(32'hbac5383c),
	.w6(32'h390cafa4),
	.w7(32'hbaab9c76),
	.w8(32'hba834206),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fe0fef),
	.w1(32'hba9df873),
	.w2(32'hbabe2ca7),
	.w3(32'hb9365e1a),
	.w4(32'hba834e7b),
	.w5(32'hbaa20bd0),
	.w6(32'hba1fd6bd),
	.w7(32'hbab95f74),
	.w8(32'hbab1c9d7),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9bf8cc),
	.w1(32'h3bc281e6),
	.w2(32'h3b9be307),
	.w3(32'h3bd44dfe),
	.w4(32'h3c13d34a),
	.w5(32'h3b6c943f),
	.w6(32'hba9e36ba),
	.w7(32'hbb12e1bc),
	.w8(32'hbbeab393),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a45dd0),
	.w1(32'hba0a8be7),
	.w2(32'hb9f26c93),
	.w3(32'hb9cf9821),
	.w4(32'hba3576b6),
	.w5(32'hba1e202a),
	.w6(32'hb9e8bffe),
	.w7(32'hba3f667f),
	.w8(32'hba11f5f5),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b838e2d),
	.w1(32'h3b8f1f62),
	.w2(32'h3b6e4c56),
	.w3(32'h3bbf3dc8),
	.w4(32'h3bc91606),
	.w5(32'h3b83e737),
	.w6(32'h3b2914bf),
	.w7(32'h3ae02c2d),
	.w8(32'hb926fad5),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99c9f4f),
	.w1(32'hba143c4c),
	.w2(32'hba0a29b9),
	.w3(32'h3a4a55b6),
	.w4(32'h3988c276),
	.w5(32'hb8ce09c8),
	.w6(32'h39edd3b6),
	.w7(32'h37bb7eb5),
	.w8(32'h39a34645),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1e5307),
	.w1(32'h3b7a6282),
	.w2(32'h3bb59233),
	.w3(32'h3b378c9f),
	.w4(32'h3b2d0a4e),
	.w5(32'h3b4cfc2c),
	.w6(32'h3afecc27),
	.w7(32'h3b151d59),
	.w8(32'h3b5c99f4),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb805be72),
	.w1(32'h3749b098),
	.w2(32'h37bda95d),
	.w3(32'hb735c652),
	.w4(32'h3816916d),
	.w5(32'h380e9be9),
	.w6(32'hb81df894),
	.w7(32'h3540d796),
	.w8(32'hb736a203),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2e0410),
	.w1(32'h3b2f142c),
	.w2(32'h3a58108d),
	.w3(32'h3ad08cf4),
	.w4(32'h39c622bc),
	.w5(32'h38d6b00a),
	.w6(32'h370ecaee),
	.w7(32'hbad37a7b),
	.w8(32'hb8bc6043),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h386242c2),
	.w1(32'h378bb6bc),
	.w2(32'h3ba7797d),
	.w3(32'h392fab31),
	.w4(32'h3ad47bee),
	.w5(32'hbaafa130),
	.w6(32'h38d82932),
	.w7(32'h3bec479f),
	.w8(32'h3907cb8a),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b463533),
	.w1(32'h3bd496bb),
	.w2(32'h3ba09191),
	.w3(32'h3bb0f52c),
	.w4(32'h3b9d0269),
	.w5(32'h3b30d4ec),
	.w6(32'h3941ff56),
	.w7(32'hb953f707),
	.w8(32'hbb0c8a71),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39adc603),
	.w1(32'h3a9a3354),
	.w2(32'hb9a0ba2e),
	.w3(32'h3b23ffac),
	.w4(32'hbacad1a8),
	.w5(32'hbb163d06),
	.w6(32'h3b1ef307),
	.w7(32'h38bb7d5e),
	.w8(32'hbb388a1e),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aacc4af),
	.w1(32'h3b618f93),
	.w2(32'hba95f5ef),
	.w3(32'h3b70f479),
	.w4(32'hbad11f86),
	.w5(32'hbae365c8),
	.w6(32'h3b2d4d62),
	.w7(32'hba85e5c5),
	.w8(32'hbb7b37d4),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e89392),
	.w1(32'h395edd84),
	.w2(32'hbaac7af2),
	.w3(32'hba717795),
	.w4(32'hbbd9561a),
	.w5(32'hbc0e870a),
	.w6(32'hbb4d6aac),
	.w7(32'h3c073176),
	.w8(32'h3b9aa797),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb04a6ed),
	.w1(32'hba6feb76),
	.w2(32'h38ff66c1),
	.w3(32'h3a273168),
	.w4(32'h3badf461),
	.w5(32'h3a88b01e),
	.w6(32'h3bf177d1),
	.w7(32'h3bb0ace0),
	.w8(32'h390b258f),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaba8053),
	.w1(32'h3ad7a40f),
	.w2(32'hbb1977be),
	.w3(32'h3b34ddb5),
	.w4(32'hbafce105),
	.w5(32'hbbb658c6),
	.w6(32'h3a1507df),
	.w7(32'hbb81e3fb),
	.w8(32'hbc265f3a),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c24db46),
	.w1(32'h3b9f4379),
	.w2(32'h3c239155),
	.w3(32'h3b8e27a3),
	.w4(32'hbac99f06),
	.w5(32'h399c6db7),
	.w6(32'h3b8421f6),
	.w7(32'h3bc53b9d),
	.w8(32'h3bc05785),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be14b45),
	.w1(32'h3c468abc),
	.w2(32'h3b34c4c2),
	.w3(32'h3a39615d),
	.w4(32'h3c4190ce),
	.w5(32'hba87a9cc),
	.w6(32'hbaeef513),
	.w7(32'h3afe104c),
	.w8(32'h3aa8ada7),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98421b8),
	.w1(32'hbb922722),
	.w2(32'hbc3658dc),
	.w3(32'h3c38c75b),
	.w4(32'h3c21382b),
	.w5(32'h3b8dc56b),
	.w6(32'h3c1f56b3),
	.w7(32'hbb96b2b6),
	.w8(32'hbc24421e),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3f3873),
	.w1(32'hbc3ec94c),
	.w2(32'hba2269da),
	.w3(32'h39c558db),
	.w4(32'hba449758),
	.w5(32'hbb9a6d83),
	.w6(32'hbbb329b9),
	.w7(32'hbbb94a12),
	.w8(32'hbbe287e1),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb06da74),
	.w1(32'hbbca06ae),
	.w2(32'hbbae3fe4),
	.w3(32'hbbdf1709),
	.w4(32'hbb5afbb7),
	.w5(32'hbc025ef5),
	.w6(32'hbc40556b),
	.w7(32'hbbc463f9),
	.w8(32'hbc244138),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc110785),
	.w1(32'h3b86919f),
	.w2(32'h37f1b9e3),
	.w3(32'h3b33bcfd),
	.w4(32'h3bb78884),
	.w5(32'h3b471695),
	.w6(32'h3b75a5d3),
	.w7(32'hb9aa3f07),
	.w8(32'hba57612a),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba14e982),
	.w1(32'h3b2fd4a2),
	.w2(32'hbc8383bc),
	.w3(32'hbb52af10),
	.w4(32'hbb772505),
	.w5(32'hbbe872ee),
	.w6(32'hbb638178),
	.w7(32'hbb44bbe4),
	.w8(32'hb90d14b7),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbde20e2),
	.w1(32'hbc2dbc27),
	.w2(32'h3b1ec1f4),
	.w3(32'hbbba518d),
	.w4(32'hbb28aba5),
	.w5(32'hbbc4baa4),
	.w6(32'hbb552a7c),
	.w7(32'hbadb742b),
	.w8(32'h3b37de0b),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3900d08e),
	.w1(32'h3b1f1bb1),
	.w2(32'h3b3c52d7),
	.w3(32'hbbe09a60),
	.w4(32'h3aca30c3),
	.w5(32'h3b36aad4),
	.w6(32'hbab0f7f3),
	.w7(32'hba905b4b),
	.w8(32'hb7aa1f1b),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3d1d9d),
	.w1(32'h3a23e58f),
	.w2(32'hbb355c92),
	.w3(32'h3acc08c5),
	.w4(32'hbbeda4be),
	.w5(32'hbbce99b3),
	.w6(32'h3ad3e309),
	.w7(32'hbc1bc2bb),
	.w8(32'hbbf722c7),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0f36a0),
	.w1(32'hba679083),
	.w2(32'h3b6131ef),
	.w3(32'h3bb0b441),
	.w4(32'h3bcd3b40),
	.w5(32'h3b34f740),
	.w6(32'hbb7387a1),
	.w7(32'h3abcbc9b),
	.w8(32'h3bfa7db2),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad00510),
	.w1(32'hbc091d1b),
	.w2(32'h3b8f2537),
	.w3(32'hbb9d8c63),
	.w4(32'hb98bddc4),
	.w5(32'h3a87eb61),
	.w6(32'hba6b162f),
	.w7(32'h39679f8b),
	.w8(32'hba9a3c6e),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad6fdde),
	.w1(32'hba52c7ae),
	.w2(32'hbbe3d724),
	.w3(32'hbb107919),
	.w4(32'h3b989d87),
	.w5(32'hbabe2b21),
	.w6(32'hbb86ba5b),
	.w7(32'hbb12b92a),
	.w8(32'hbb41485b),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7a1260),
	.w1(32'h3c29d8f8),
	.w2(32'h3bd0231d),
	.w3(32'h3b9d1466),
	.w4(32'hbb796412),
	.w5(32'h39facc14),
	.w6(32'h3ad9749c),
	.w7(32'hbc20d953),
	.w8(32'hbc5127c0),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e85767),
	.w1(32'hbb5ecef5),
	.w2(32'hbb13ea86),
	.w3(32'h3bcac99c),
	.w4(32'hbb8f68a9),
	.w5(32'hbc3d8dab),
	.w6(32'hbb2d0288),
	.w7(32'h3be9aa81),
	.w8(32'h3bce89ea),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf87029),
	.w1(32'hbc155371),
	.w2(32'h3a9f0288),
	.w3(32'hbc196259),
	.w4(32'h3af7a887),
	.w5(32'hbb30884f),
	.w6(32'h3bd50f89),
	.w7(32'h3b975326),
	.w8(32'hb9c3d437),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5e04b8),
	.w1(32'hbbc3ab28),
	.w2(32'hbca7afff),
	.w3(32'hbb2cf318),
	.w4(32'hbc7fdb80),
	.w5(32'hbcad1518),
	.w6(32'hbb810ef6),
	.w7(32'hbcf4bd91),
	.w8(32'hbd0060a9),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc05556),
	.w1(32'hbcadb0f0),
	.w2(32'hb9990f45),
	.w3(32'hbcf39737),
	.w4(32'h3bb6bbda),
	.w5(32'h3b2fc4b5),
	.w6(32'hbd08b46d),
	.w7(32'hbbc84c15),
	.w8(32'hbb828d1e),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f12436),
	.w1(32'h3a7abbff),
	.w2(32'h3b144b5b),
	.w3(32'h3baa95a9),
	.w4(32'h3b36c673),
	.w5(32'h3ba44c64),
	.w6(32'hbb44574f),
	.w7(32'hbbbf4d93),
	.w8(32'hbb21c8d0),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bdce99),
	.w1(32'h3a40587b),
	.w2(32'hbb82ba59),
	.w3(32'hba9262ce),
	.w4(32'hbc1045d9),
	.w5(32'hbbf799bc),
	.w6(32'hbb7a0b2f),
	.w7(32'hbc069b81),
	.w8(32'hbb20e724),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb45b6e0),
	.w1(32'hbbadc955),
	.w2(32'h3c4c4993),
	.w3(32'hbaeebd50),
	.w4(32'hba484512),
	.w5(32'h391f40eb),
	.w6(32'h3b3ae519),
	.w7(32'hbb055e03),
	.w8(32'hbbed06d5),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd6bf59),
	.w1(32'hba974b87),
	.w2(32'hbb23b1ee),
	.w3(32'h3af54606),
	.w4(32'hbba02be9),
	.w5(32'hbbd5d827),
	.w6(32'hbb91a6cc),
	.w7(32'h38e7cbe6),
	.w8(32'hbb384718),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba674ec5),
	.w1(32'h3a3ed36f),
	.w2(32'hbbe964e0),
	.w3(32'h3a8dc508),
	.w4(32'h3c4eef78),
	.w5(32'h3b868128),
	.w6(32'hb9e313fa),
	.w7(32'hbb715779),
	.w8(32'hbbfe8dd6),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2b0ef7),
	.w1(32'h3c1bc9a5),
	.w2(32'h3c3beb48),
	.w3(32'h3b3ca786),
	.w4(32'hba619c26),
	.w5(32'hbb6263fb),
	.w6(32'hbc10ea45),
	.w7(32'hbc02fdc3),
	.w8(32'hbbe9dec7),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7db912),
	.w1(32'hbbbaa33a),
	.w2(32'h3be70c46),
	.w3(32'hbb0fb5a4),
	.w4(32'h3b5db87c),
	.w5(32'hbac2665f),
	.w6(32'hbbb9f2a2),
	.w7(32'h3bf9c822),
	.w8(32'hbb2ca989),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba443b9b),
	.w1(32'h3a807032),
	.w2(32'hba8d72f6),
	.w3(32'h3a9b0ed2),
	.w4(32'hbc0cdc3e),
	.w5(32'hbbbd7ed6),
	.w6(32'hb9c45f8e),
	.w7(32'hbb33adc9),
	.w8(32'hb9e65e41),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbb56b8),
	.w1(32'hbb2da27f),
	.w2(32'h3c074c89),
	.w3(32'hb9c4f880),
	.w4(32'h3c8a4e5a),
	.w5(32'h3c02e69a),
	.w6(32'hbb7f4384),
	.w7(32'hbbb89d55),
	.w8(32'hbc2cedd2),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1e09e9),
	.w1(32'h3c191c22),
	.w2(32'h3c2b7321),
	.w3(32'h391e3fc0),
	.w4(32'hbc16cb6d),
	.w5(32'hbb2d9ec5),
	.w6(32'hbb8d445d),
	.w7(32'hbaa799e9),
	.w8(32'h3a25231d),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c488da0),
	.w1(32'h3b166598),
	.w2(32'h3b9b2108),
	.w3(32'h3b295f32),
	.w4(32'hb99527f8),
	.w5(32'hba8cc98e),
	.w6(32'hba5ab777),
	.w7(32'hbb37a6c3),
	.w8(32'hbbb1cdd6),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb872f92),
	.w1(32'hbbbcf16f),
	.w2(32'h37229226),
	.w3(32'hbb7bced4),
	.w4(32'hbb94b0c2),
	.w5(32'hba45125f),
	.w6(32'hbbc5a53c),
	.w7(32'h3b92442d),
	.w8(32'h3bd6e19e),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3c7f4a),
	.w1(32'hbb0ab684),
	.w2(32'hbbbde9bb),
	.w3(32'hba802312),
	.w4(32'hbb05f4f0),
	.w5(32'hbbf0fb9b),
	.w6(32'h39c7747f),
	.w7(32'hbc0ad056),
	.w8(32'hbc830333),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc22fa08),
	.w1(32'hbb88ee00),
	.w2(32'hbc254b5f),
	.w3(32'hbb938dd0),
	.w4(32'h3b54fc74),
	.w5(32'h3a4b4c2d),
	.w6(32'hbc35ecc8),
	.w7(32'h3b8cd831),
	.w8(32'h3b1c7dca),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ce2be),
	.w1(32'h3c421360),
	.w2(32'h3c200d59),
	.w3(32'hbc03c503),
	.w4(32'h3c103ead),
	.w5(32'h3c7d838e),
	.w6(32'h3b3a053f),
	.w7(32'h3d0c0ba0),
	.w8(32'h3d523a72),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c51d636),
	.w1(32'h3bda19a9),
	.w2(32'hbbed6ae1),
	.w3(32'h3c8343d1),
	.w4(32'hbb32c953),
	.w5(32'h3b3a284e),
	.w6(32'h3d2a52b4),
	.w7(32'hbc32a340),
	.w8(32'hbbc0743d),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb103619),
	.w1(32'h3a085d75),
	.w2(32'h3bc911af),
	.w3(32'h3b3f05ba),
	.w4(32'h3ae479b5),
	.w5(32'hb9fce44f),
	.w6(32'hbb414ae6),
	.w7(32'h3b697948),
	.w8(32'hbaa4534c),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39818076),
	.w1(32'h3ac925c3),
	.w2(32'h3c2098a5),
	.w3(32'h3ab147af),
	.w4(32'hbb249907),
	.w5(32'hbb356a54),
	.w6(32'h38170cf4),
	.w7(32'h3b0dfc79),
	.w8(32'h3a2f660d),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1e8a97),
	.w1(32'h3b99e099),
	.w2(32'h3a09a365),
	.w3(32'hbadcff5a),
	.w4(32'h3a37b17f),
	.w5(32'hbb81c318),
	.w6(32'h3b505a9c),
	.w7(32'h3abf2c78),
	.w8(32'hbc090e90),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb98a96a),
	.w1(32'hba47b92d),
	.w2(32'h3b2d5a6f),
	.w3(32'h3b15d9da),
	.w4(32'hb9944671),
	.w5(32'hbb8314c4),
	.w6(32'hbb1bf80b),
	.w7(32'hbbfe5a30),
	.w8(32'hbc327d3a),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be55554),
	.w1(32'h3c085d95),
	.w2(32'h3c28fcc6),
	.w3(32'hba96b60f),
	.w4(32'h3c808770),
	.w5(32'h3b90e435),
	.w6(32'hbb802e38),
	.w7(32'h3c55bc29),
	.w8(32'h3bbba185),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0c872b),
	.w1(32'h3ad9201c),
	.w2(32'h3bbcafec),
	.w3(32'hbc08339c),
	.w4(32'h3aaa8cee),
	.w5(32'hbaa8d0a3),
	.w6(32'hbb9d0ed9),
	.w7(32'h3bdbc309),
	.w8(32'hba00be1d),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa90417),
	.w1(32'hb7384eca),
	.w2(32'hbb3491f4),
	.w3(32'hb890bc6f),
	.w4(32'hbc0be387),
	.w5(32'hbb26a591),
	.w6(32'hb9da39e3),
	.w7(32'hbc1d6e12),
	.w8(32'hbb0a8884),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaab535a),
	.w1(32'hbaa1ddc2),
	.w2(32'hbbace311),
	.w3(32'h3b875bf3),
	.w4(32'h3c642a64),
	.w5(32'h3b7be7e5),
	.w6(32'h3bd08b74),
	.w7(32'hbbde3740),
	.w8(32'hbc0e8280),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb0572d),
	.w1(32'hba451a01),
	.w2(32'hbb5b3e70),
	.w3(32'hba65871e),
	.w4(32'hbadfe47e),
	.w5(32'hbb5b0e88),
	.w6(32'hbc128ce5),
	.w7(32'hbbfeeb2b),
	.w8(32'hbc4ddcf4),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4d9cb4),
	.w1(32'h3b15ae09),
	.w2(32'h3ab8529a),
	.w3(32'h3a6ff247),
	.w4(32'hbb1ddd23),
	.w5(32'hbb9442d9),
	.w6(32'hbba7aab8),
	.w7(32'hbb0e51f5),
	.w8(32'hbb95c608),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb26421f),
	.w1(32'h38314fba),
	.w2(32'h3a04c608),
	.w3(32'h39fba2f9),
	.w4(32'hba97f831),
	.w5(32'hbb18ad30),
	.w6(32'h3ae2f1fe),
	.w7(32'hb9ec43fa),
	.w8(32'hbb334318),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule