module layer_6_featuremap_122(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 2048;
	parameter IMG_SIZE = 52;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b499c42),
	.w1(32'hb9f673b4),
	.w2(32'h3b95a5dd),
	.w3(32'hbc12e44c),
	.w4(32'hbb14a844),
	.w5(32'hbb879b55),
	.w6(32'h3b2d12d2),
	.w7(32'h3b330ab6),
	.w8(32'h3b1c0e2a),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaca5de),
	.w1(32'hb9728dd5),
	.w2(32'hbb2859b4),
	.w3(32'hbb764680),
	.w4(32'hbbea4e5c),
	.w5(32'hbbb4b462),
	.w6(32'h3b8a5a65),
	.w7(32'h3bdf2782),
	.w8(32'h3b87b93c),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ddb8e9),
	.w1(32'h3c03e54f),
	.w2(32'hbb8caf30),
	.w3(32'hbb1f8480),
	.w4(32'hbc0d3983),
	.w5(32'h3c0b4291),
	.w6(32'h3c417930),
	.w7(32'h3b19019a),
	.w8(32'hb99d6524),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c10fba7),
	.w1(32'h3b449786),
	.w2(32'h3b58740f),
	.w3(32'h3b2c3985),
	.w4(32'h3b42f61c),
	.w5(32'h3b22aa5f),
	.w6(32'h3b4af2f3),
	.w7(32'h3aea7d98),
	.w8(32'h3bbb9587),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacd618b),
	.w1(32'h3ce18cd6),
	.w2(32'hbd5abb53),
	.w3(32'h3cbb503c),
	.w4(32'hbcfa106a),
	.w5(32'h3c244deb),
	.w6(32'hbd1ba2c6),
	.w7(32'h3d611684),
	.w8(32'hbd4ec605),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4b13cc),
	.w1(32'hba98bdaf),
	.w2(32'hbb8c1d28),
	.w3(32'hbbecea5c),
	.w4(32'h3a3428b8),
	.w5(32'hba490350),
	.w6(32'hbb4d9711),
	.w7(32'hbaf80d90),
	.w8(32'h3acf70cd),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a2e2b),
	.w1(32'hbc0b72e7),
	.w2(32'h3aad937f),
	.w3(32'hbc4a25e9),
	.w4(32'hbc30556d),
	.w5(32'hbbec60a2),
	.w6(32'hbbed0e10),
	.w7(32'hbac5ea35),
	.w8(32'hbb340a4c),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae59730),
	.w1(32'h3be5de54),
	.w2(32'hbc138772),
	.w3(32'h39f30f67),
	.w4(32'hbc91bdc2),
	.w5(32'h3c0ba8b2),
	.w6(32'hbc9922b9),
	.w7(32'h3cc11b30),
	.w8(32'hbc9be3d4),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5161c6),
	.w1(32'h3d5ae8eb),
	.w2(32'hbd847377),
	.w3(32'h3d0ba912),
	.w4(32'hbd79dd7e),
	.w5(32'h3cc27a13),
	.w6(32'hbdb38192),
	.w7(32'h3dc17eeb),
	.w8(32'hbd4392a2),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c359e44),
	.w1(32'hbb16fcee),
	.w2(32'h3b4fbd22),
	.w3(32'hbbaac000),
	.w4(32'h3aa0e014),
	.w5(32'h3b06daf0),
	.w6(32'h3a7065ca),
	.w7(32'hb90e09af),
	.w8(32'h3b8bba9c),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9f3444),
	.w1(32'h3b38b2ea),
	.w2(32'hb826eaf1),
	.w3(32'h3bc7b1d4),
	.w4(32'hbb91aa33),
	.w5(32'hbb564856),
	.w6(32'hbb90b600),
	.w7(32'h3b3ec9bb),
	.w8(32'hbbf12183),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c25ec61),
	.w1(32'h3c309098),
	.w2(32'hbabde40a),
	.w3(32'hbae07276),
	.w4(32'h3b13497f),
	.w5(32'h3c1441b1),
	.w6(32'h3bac8c88),
	.w7(32'hbb73aa24),
	.w8(32'h3aa66806),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5a83cd),
	.w1(32'hb9a3ee5f),
	.w2(32'h3a6b8d94),
	.w3(32'hbb7bca0e),
	.w4(32'h39681f2f),
	.w5(32'hba215ff4),
	.w6(32'h3af3f1ce),
	.w7(32'h3abd0667),
	.w8(32'h3afe7f12),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3828837d),
	.w1(32'h3cc87e6b),
	.w2(32'hbd5ec241),
	.w3(32'hbcb868dc),
	.w4(32'h3d0fea5e),
	.w5(32'hbc11cb8c),
	.w6(32'hbbf635b7),
	.w7(32'h3d41d042),
	.w8(32'hbc85445a),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d2e06bb),
	.w1(32'h3b604a96),
	.w2(32'hba3ea4a6),
	.w3(32'h39561662),
	.w4(32'h3b7c41f3),
	.w5(32'h3b22cec4),
	.w6(32'hbbd89242),
	.w7(32'hbb04a66f),
	.w8(32'h3b109d73),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3bc487),
	.w1(32'hbbb002c0),
	.w2(32'h381520a2),
	.w3(32'hb8fc5434),
	.w4(32'hbae14b92),
	.w5(32'hbb9141f6),
	.w6(32'hbab48629),
	.w7(32'hbbbdacfb),
	.w8(32'hb98f4750),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b902320),
	.w1(32'hbbae47c2),
	.w2(32'hbc4e0f3b),
	.w3(32'h39511cdb),
	.w4(32'hbbbe5136),
	.w5(32'hbc93fae2),
	.w6(32'hbc4ec98f),
	.w7(32'hbce80ad9),
	.w8(32'hbc127782),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc83e451),
	.w1(32'hbb7ef63e),
	.w2(32'h3bf8ab46),
	.w3(32'h39d0cc3d),
	.w4(32'h3b661617),
	.w5(32'hb79028ec),
	.w6(32'h3b232921),
	.w7(32'h3acc0e45),
	.w8(32'h3bfc8cce),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb976d744),
	.w1(32'hbba63d10),
	.w2(32'hbb5a8000),
	.w3(32'hba166f5c),
	.w4(32'h3abb90b6),
	.w5(32'h3b082dad),
	.w6(32'hbb1887b8),
	.w7(32'hbaf987dc),
	.w8(32'hbb3b5c2e),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaab5850),
	.w1(32'hbb5a5a17),
	.w2(32'h3bb8bb1a),
	.w3(32'h3a6ee550),
	.w4(32'hb851f1bc),
	.w5(32'h3b54e77b),
	.w6(32'hbbaa91f5),
	.w7(32'h3bd8c076),
	.w8(32'hbba4ed67),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a62e22e),
	.w1(32'h3a05f759),
	.w2(32'h3a8db6c5),
	.w3(32'h39fb6cc8),
	.w4(32'hbb2611a3),
	.w5(32'hbb1605b8),
	.w6(32'hb9ab6f15),
	.w7(32'hbb024cd0),
	.w8(32'h3a3d1c81),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcd0015),
	.w1(32'h3baefc11),
	.w2(32'h3bdfedeb),
	.w3(32'h3b902b94),
	.w4(32'h3bb4d5d6),
	.w5(32'h3bbf211e),
	.w6(32'h3c0fd948),
	.w7(32'h3b615a30),
	.w8(32'h3c201602),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2a0f95),
	.w1(32'hbb0a0d0c),
	.w2(32'hbb8efdf0),
	.w3(32'hbcc485df),
	.w4(32'hbbb8f60b),
	.w5(32'h3b8059af),
	.w6(32'hbb3f28e8),
	.w7(32'hbc8b0919),
	.w8(32'h3b1d260c),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb085fca),
	.w1(32'h3c00d187),
	.w2(32'h3b81b41c),
	.w3(32'hbc98b698),
	.w4(32'h3cf63899),
	.w5(32'hbb5ca086),
	.w6(32'hbb1c9848),
	.w7(32'hbcdd1a7c),
	.w8(32'h3ab42969),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae70e41),
	.w1(32'hbaad3e9e),
	.w2(32'h3bb2d6b2),
	.w3(32'hbc03bf11),
	.w4(32'h3c5c6e7e),
	.w5(32'hbac0a63a),
	.w6(32'h3a20471d),
	.w7(32'hbba9b39f),
	.w8(32'h3c4cd93d),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd36b6d),
	.w1(32'h3ca1b62e),
	.w2(32'h3b628c7b),
	.w3(32'h3c0b9d32),
	.w4(32'h3c4505a7),
	.w5(32'h3c05ba56),
	.w6(32'h3b335671),
	.w7(32'h3b41b4b6),
	.w8(32'h3c24fbf6),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af3dee1),
	.w1(32'h3b64744c),
	.w2(32'h3c3fad39),
	.w3(32'h3c02d227),
	.w4(32'h3be29d31),
	.w5(32'h3bdd4937),
	.w6(32'h3c151d36),
	.w7(32'h3b313671),
	.w8(32'h3c3c81d0),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8e6570),
	.w1(32'hbb1b5535),
	.w2(32'hba141f1d),
	.w3(32'hb9aca328),
	.w4(32'h3993e1c3),
	.w5(32'hb918fb1f),
	.w6(32'hbaeb4dc1),
	.w7(32'h39bd94f2),
	.w8(32'hba3566e5),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4a7e0d),
	.w1(32'hbb1a8b53),
	.w2(32'hb9276f53),
	.w3(32'h3a08a4dd),
	.w4(32'hbad4c7d7),
	.w5(32'hbb1d587d),
	.w6(32'hba8da79b),
	.w7(32'hb8f4f781),
	.w8(32'hbb46b371),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aac1ae1),
	.w1(32'hbd288c97),
	.w2(32'h3d9d117d),
	.w3(32'h3cf076ac),
	.w4(32'hbc93c8df),
	.w5(32'h3d4a4d60),
	.w6(32'h3d6d7fa4),
	.w7(32'h3d418a72),
	.w8(32'h3ca95ab1),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be5e68f),
	.w1(32'h3cd0966c),
	.w2(32'hbb9fb9a9),
	.w3(32'h3cd64592),
	.w4(32'hbc8fad79),
	.w5(32'hbb615106),
	.w6(32'hbd15c060),
	.w7(32'h3cd2de72),
	.w8(32'hbca96b62),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbae9a4d),
	.w1(32'h3bad6434),
	.w2(32'h3c1ca61a),
	.w3(32'h3b426fda),
	.w4(32'h39450a00),
	.w5(32'h3b22da52),
	.w6(32'hbb3105d7),
	.w7(32'h3a93a2db),
	.w8(32'h3c1c191a),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba52cd9f),
	.w1(32'hbc9cbf96),
	.w2(32'h3c43858d),
	.w3(32'hbb357192),
	.w4(32'hbb5883f4),
	.w5(32'hbb0b26e6),
	.w6(32'hbb7e5610),
	.w7(32'hbcab0c94),
	.w8(32'h3c6ab1f6),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6f47ba),
	.w1(32'h3d3e3c30),
	.w2(32'h3cb03e8c),
	.w3(32'h3c9d5ce9),
	.w4(32'h3d8210ee),
	.w5(32'hbc4a29c8),
	.w6(32'h3ccaa135),
	.w7(32'h3d96cc12),
	.w8(32'h3d021bd5),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d3dd13c),
	.w1(32'h3b3651db),
	.w2(32'hbab59934),
	.w3(32'hbb20e4c1),
	.w4(32'hba28139b),
	.w5(32'h3ac34d45),
	.w6(32'h3a9964ee),
	.w7(32'hb977775b),
	.w8(32'h3b01aff0),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc1406c),
	.w1(32'h3b92b290),
	.w2(32'h3b87b8b4),
	.w3(32'h3bc31c31),
	.w4(32'h3b4e47c7),
	.w5(32'hbac44d9e),
	.w6(32'h3ae82474),
	.w7(32'hbab1baae),
	.w8(32'h39d76385),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4a30fd),
	.w1(32'h3ba40b55),
	.w2(32'hbb7eafa7),
	.w3(32'hbb87b025),
	.w4(32'h3b44d42f),
	.w5(32'hba4cc03f),
	.w6(32'hbb02e927),
	.w7(32'h390cb068),
	.w8(32'hbac10982),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afa37c5),
	.w1(32'h3b663419),
	.w2(32'h3b803a81),
	.w3(32'h3b26f823),
	.w4(32'h3b20a322),
	.w5(32'hba7f8904),
	.w6(32'h3b576e41),
	.w7(32'h3b0f9ebd),
	.w8(32'h388263b5),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a99dbce),
	.w1(32'hbb8c09dd),
	.w2(32'hbbd753f0),
	.w3(32'h3a175ada),
	.w4(32'hbb283647),
	.w5(32'h3c117839),
	.w6(32'hbc95ff97),
	.w7(32'hbb9f5e75),
	.w8(32'h3c62e449),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8a006a),
	.w1(32'h3d155dd9),
	.w2(32'hbc6897ed),
	.w3(32'h3d243d35),
	.w4(32'hbd282380),
	.w5(32'h3cff7237),
	.w6(32'hbd55423d),
	.w7(32'h3d8e2edd),
	.w8(32'hbc66b351),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc36fca1),
	.w1(32'hbbbf96a5),
	.w2(32'hbc582f51),
	.w3(32'h3c063f87),
	.w4(32'hbc804b70),
	.w5(32'h3c0ffe2a),
	.w6(32'hbbd94113),
	.w7(32'h3d000070),
	.w8(32'hbaa327f2),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0e5124),
	.w1(32'hbaca5e65),
	.w2(32'h39ada67e),
	.w3(32'h3916d4fb),
	.w4(32'h3944e6c3),
	.w5(32'hbb302ad5),
	.w6(32'h3aa9b3db),
	.w7(32'hbaa211b9),
	.w8(32'h3a70f928),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb168efd),
	.w1(32'h3bcbeb53),
	.w2(32'h3be3b34b),
	.w3(32'h3af3dbf9),
	.w4(32'h3ba68c36),
	.w5(32'h3c5c46ed),
	.w6(32'h3b7229be),
	.w7(32'h3be3059c),
	.w8(32'h3c447c47),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c439314),
	.w1(32'h3c4ed6d0),
	.w2(32'h3acff0fe),
	.w3(32'h3c0fcac4),
	.w4(32'h3bab6d9d),
	.w5(32'h3bae2c8e),
	.w6(32'h3b024981),
	.w7(32'h3bd5525d),
	.w8(32'h3b753122),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeb1c64),
	.w1(32'hbaef5338),
	.w2(32'h3b3a62c2),
	.w3(32'hbb04e062),
	.w4(32'hbab8fac0),
	.w5(32'h3b18854a),
	.w6(32'h3acc6d8a),
	.w7(32'hba90d73c),
	.w8(32'h3b132cc3),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0d727f),
	.w1(32'hbccda601),
	.w2(32'h3a4672f7),
	.w3(32'hbcc2e5ec),
	.w4(32'hbc958a54),
	.w5(32'hbbba43cb),
	.w6(32'hbb8c86f8),
	.w7(32'hbc8fbd35),
	.w8(32'hbbd9240f),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7a12df),
	.w1(32'h3b7afe87),
	.w2(32'h3c3b755a),
	.w3(32'hbb85423e),
	.w4(32'hbbd097cb),
	.w5(32'hbb5e0b0f),
	.w6(32'h3addaac4),
	.w7(32'h3be1afbd),
	.w8(32'h3bf26048),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c45a064),
	.w1(32'h3b9752c5),
	.w2(32'hbbaa6442),
	.w3(32'hbbaf3d7e),
	.w4(32'h3a8586ae),
	.w5(32'h3a6533b5),
	.w6(32'hbc5b7d6a),
	.w7(32'hbc84b0c4),
	.w8(32'h3bbfad0e),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4a8c33),
	.w1(32'h3ba0e3ce),
	.w2(32'h3b815126),
	.w3(32'h3a2d2d2d),
	.w4(32'h39aa9888),
	.w5(32'h3bb10195),
	.w6(32'h3a98db99),
	.w7(32'h3a6779d3),
	.w8(32'h3afb7696),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8cda61),
	.w1(32'hbd19f918),
	.w2(32'h3d130ad0),
	.w3(32'hbd073425),
	.w4(32'h3d14ed05),
	.w5(32'hbc6b35bc),
	.w6(32'h3d4638c5),
	.w7(32'hbdb016c6),
	.w8(32'h3d00b4b6),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c68a37f),
	.w1(32'hba3ffebf),
	.w2(32'h3b4fc0ed),
	.w3(32'hbab0e0e7),
	.w4(32'h3b2fa410),
	.w5(32'hbb69ecc5),
	.w6(32'h3b95d3b3),
	.w7(32'h3a8ebf59),
	.w8(32'h3b99b709),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba28bdf),
	.w1(32'h3b899e17),
	.w2(32'h3b05e749),
	.w3(32'hbbae73d5),
	.w4(32'hbbc5c4a3),
	.w5(32'hba00a03c),
	.w6(32'hba924ff4),
	.w7(32'hbb5652ef),
	.w8(32'h3b1f779e),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9c6944),
	.w1(32'hb6df2d10),
	.w2(32'hb9c6d921),
	.w3(32'hbaa7eaec),
	.w4(32'hbb0ec67e),
	.w5(32'hb9872cd2),
	.w6(32'hbadafeaa),
	.w7(32'hbaa77157),
	.w8(32'h3ae4604f),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3b4ec5),
	.w1(32'h3c1747c6),
	.w2(32'h3bfe1016),
	.w3(32'hbb78edca),
	.w4(32'hbb11e65c),
	.w5(32'hbb89e658),
	.w6(32'h3c01a622),
	.w7(32'h3bf5ce4a),
	.w8(32'h3c13dfd8),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c287a60),
	.w1(32'h3b313b5a),
	.w2(32'h3b394558),
	.w3(32'hbb71034e),
	.w4(32'hbb22b212),
	.w5(32'hbb46d996),
	.w6(32'h3bcd9ca6),
	.w7(32'h3b1e3b57),
	.w8(32'h3bedf3c0),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba1cd8d),
	.w1(32'hbbe881b2),
	.w2(32'h3a67eab5),
	.w3(32'h3a90c428),
	.w4(32'h3b40bd33),
	.w5(32'hbb238605),
	.w6(32'hbb97bf96),
	.w7(32'hbbc2130a),
	.w8(32'hbaaa6f15),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7752eea),
	.w1(32'hb9e5cd2c),
	.w2(32'h3b87f75d),
	.w3(32'hbb87fba9),
	.w4(32'h3a71d6fe),
	.w5(32'hbb27611c),
	.w6(32'h3a7193f8),
	.w7(32'h3bda9961),
	.w8(32'h3ae304fe),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad5d6cb),
	.w1(32'h3ad64578),
	.w2(32'h3b67dd8e),
	.w3(32'h3bc881ed),
	.w4(32'h3c5e9eba),
	.w5(32'h3b58bbf0),
	.w6(32'h3bf57821),
	.w7(32'h3c801eb8),
	.w8(32'h3c322d98),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b36090e),
	.w1(32'h3b089ac1),
	.w2(32'h3b301d65),
	.w3(32'h3b26b1cf),
	.w4(32'h3b4ca4cc),
	.w5(32'h3b1b43ff),
	.w6(32'h3b82830a),
	.w7(32'h3b9b8530),
	.w8(32'h3b6253a2),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b879091),
	.w1(32'h3bc95c42),
	.w2(32'h3b7346d4),
	.w3(32'h3b7e990e),
	.w4(32'h3c1350df),
	.w5(32'h3bcf40a5),
	.w6(32'hbb90e5eb),
	.w7(32'hbb88edeb),
	.w8(32'h3ba036ed),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbc8fe7),
	.w1(32'hbb937b8d),
	.w2(32'hba91a3ad),
	.w3(32'hbbc1bb8a),
	.w4(32'hbb02ea6a),
	.w5(32'hbbaa1f30),
	.w6(32'h39ce3941),
	.w7(32'h3b43e25b),
	.w8(32'h39f57c5a),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8808d7),
	.w1(32'h3b38c0b0),
	.w2(32'h3b999847),
	.w3(32'h3bb4c77c),
	.w4(32'h3c4772a7),
	.w5(32'h3c4bf036),
	.w6(32'h3bd9b2b5),
	.w7(32'h3c57961c),
	.w8(32'h3c129330),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d7f1f1),
	.w1(32'h3b6172e3),
	.w2(32'hbc112f33),
	.w3(32'h3bb2970e),
	.w4(32'h3bd15ac2),
	.w5(32'h3b32a705),
	.w6(32'h3c245bcc),
	.w7(32'h3b1b80e9),
	.w8(32'h3c1cc41f),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabe1893),
	.w1(32'h3c43738c),
	.w2(32'h3c6dad36),
	.w3(32'h3c818227),
	.w4(32'h3c92199b),
	.w5(32'h3c468e01),
	.w6(32'h3c907dfc),
	.w7(32'h3cb471a5),
	.w8(32'h3c425a00),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

endmodule