module layer_10_featuremap_219(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h34123ed4),
	.w1(32'hb4a2feba),
	.w2(32'h3588d0ee),
	.w3(32'hb44e2c8f),
	.w4(32'h34bbb713),
	.w5(32'h358357c3),
	.w6(32'hb55ed86c),
	.w7(32'hb5639141),
	.w8(32'h334dbdca),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb69e45aa),
	.w1(32'hb7254623),
	.w2(32'h35d2ca2c),
	.w3(32'hb7647cb7),
	.w4(32'hb7640027),
	.w5(32'h340c9e53),
	.w6(32'hb6be1c32),
	.w7(32'hb6d0aead),
	.w8(32'h36a40d0d),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb43804c9),
	.w1(32'hb5d85539),
	.w2(32'hb5b3eded),
	.w3(32'h34bf477e),
	.w4(32'hb5241e5c),
	.w5(32'hb507df9f),
	.w6(32'hb41636ef),
	.w7(32'hb54089bc),
	.w8(32'hb5a6e61d),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb621696b),
	.w1(32'hb520f548),
	.w2(32'h362405ea),
	.w3(32'hb639a16a),
	.w4(32'h347c2d89),
	.w5(32'h361cec90),
	.w6(32'hb64588fc),
	.w7(32'h35d51b53),
	.w8(32'h3557e10b),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3644b03e),
	.w1(32'h36770d6f),
	.w2(32'h3698ab73),
	.w3(32'h35f8b18d),
	.w4(32'h35d0f5c8),
	.w5(32'h36219cb8),
	.w6(32'h33a05be1),
	.w7(32'h35cf117c),
	.w8(32'hb5e384e8),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5ae2af3),
	.w1(32'h34a3a471),
	.w2(32'hb4a636a6),
	.w3(32'hb6003d2b),
	.w4(32'h32d812a5),
	.w5(32'hb5b5cb21),
	.w6(32'hb5187336),
	.w7(32'hb4985514),
	.w8(32'hb2d71ed9),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6925ead),
	.w1(32'hb63b0c95),
	.w2(32'hb6bc60a4),
	.w3(32'h364429fd),
	.w4(32'h36b93cea),
	.w5(32'hb7421701),
	.w6(32'h36266ca8),
	.w7(32'h3666299e),
	.w8(32'hb772f984),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37c8713f),
	.w1(32'h379523c0),
	.w2(32'h380afd76),
	.w3(32'h37bd1715),
	.w4(32'h37e2e357),
	.w5(32'h380200d4),
	.w6(32'h37232761),
	.w7(32'h37f216f6),
	.w8(32'h38255a0c),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb4988eec),
	.w1(32'h36296e0a),
	.w2(32'h3802084c),
	.w3(32'hb581ef34),
	.w4(32'h3606fd46),
	.w5(32'h3803715e),
	.w6(32'h365ca397),
	.w7(32'h3719890c),
	.w8(32'h3817a059),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb677c91f),
	.w1(32'hb7fd551f),
	.w2(32'h3825aa50),
	.w3(32'hb80c6f3c),
	.w4(32'hb81bc959),
	.w5(32'h381c4be8),
	.w6(32'hb6f613e6),
	.w7(32'hb7c8e181),
	.w8(32'h38181788),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3816b614),
	.w1(32'h37910056),
	.w2(32'h378488cc),
	.w3(32'h37a6a742),
	.w4(32'h3794a6c2),
	.w5(32'h3743e82c),
	.w6(32'h3780edfc),
	.w7(32'h37340702),
	.w8(32'hb68cef62),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h380277d7),
	.w1(32'h37238608),
	.w2(32'hb773b78c),
	.w3(32'h37bca251),
	.w4(32'h36eb2f2c),
	.w5(32'hb7dfaf5d),
	.w6(32'h38178db0),
	.w7(32'h372d0096),
	.w8(32'hb7ac5339),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6338372),
	.w1(32'hb7cfd27e),
	.w2(32'h381fe245),
	.w3(32'hb72fe728),
	.w4(32'hb74b6d0f),
	.w5(32'h38394905),
	.w6(32'hb79a3f46),
	.w7(32'hb67a9b03),
	.w8(32'h383c0a8b),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h369fd58c),
	.w1(32'h36e06e20),
	.w2(32'h377b65f3),
	.w3(32'h3740e925),
	.w4(32'h36bbdbc7),
	.w5(32'h37945dfd),
	.w6(32'h35eca530),
	.w7(32'h36eaab17),
	.w8(32'h377d401d),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7630e17),
	.w1(32'hb7a4c38f),
	.w2(32'h37810559),
	.w3(32'hb64c0a8e),
	.w4(32'hb796201a),
	.w5(32'h375c2416),
	.w6(32'h3642b0f3),
	.w7(32'hb3e03ad1),
	.w8(32'h37a265fd),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7b33113),
	.w1(32'hb7c04dcf),
	.w2(32'h37db83d7),
	.w3(32'hb76815be),
	.w4(32'h36bbf181),
	.w5(32'h385838ae),
	.w6(32'h361c1e0b),
	.w7(32'h37184a71),
	.w8(32'h3876371e),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36f6fdac),
	.w1(32'h349b4845),
	.w2(32'hb6dbb5b0),
	.w3(32'hb7956631),
	.w4(32'hb81262b9),
	.w5(32'hb790815a),
	.w6(32'h3761032c),
	.w7(32'hb695d331),
	.w8(32'hb68f5346),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5bd5057),
	.w1(32'hb6a57541),
	.w2(32'h3810488e),
	.w3(32'hb434f77d),
	.w4(32'h3730d06d),
	.w5(32'h37ef36ec),
	.w6(32'h34c5eea2),
	.w7(32'h360f3b99),
	.w8(32'h37935899),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb773ae76),
	.w1(32'hb67c4029),
	.w2(32'h381dcccf),
	.w3(32'hb6cabf7a),
	.w4(32'h378047e8),
	.w5(32'h384dd2c1),
	.w6(32'hb5ffc22f),
	.w7(32'h379594f7),
	.w8(32'h38253f86),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h347d0209),
	.w1(32'h34549b2d),
	.w2(32'hb4379f77),
	.w3(32'h33357835),
	.w4(32'h3515a558),
	.w5(32'h33b454ae),
	.w6(32'hb58307f5),
	.w7(32'hb4f4d80d),
	.w8(32'hb4a52607),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb3f77163),
	.w1(32'h3504b9fe),
	.w2(32'hb562af14),
	.w3(32'h34c2c59a),
	.w4(32'h34ec81ed),
	.w5(32'hb536e35b),
	.w6(32'hb60894cc),
	.w7(32'hb59ab3c9),
	.w8(32'hb5537d80),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3578ec2e),
	.w1(32'h36e41582),
	.w2(32'h376fb165),
	.w3(32'hb6a12727),
	.w4(32'h35bbb7bb),
	.w5(32'h36eede30),
	.w6(32'h3723c6e7),
	.w7(32'h36f16a1c),
	.w8(32'h371a3a1b),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb82d3981),
	.w1(32'hb86dc75b),
	.w2(32'h38801d2e),
	.w3(32'h36561af7),
	.w4(32'hb6981098),
	.w5(32'h389cea68),
	.w6(32'h38a423cf),
	.w7(32'h38620562),
	.w8(32'h390c7de8),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb80239e3),
	.w1(32'hb8385f57),
	.w2(32'h38001115),
	.w3(32'hb8455736),
	.w4(32'hb82dfac9),
	.w5(32'h384041e3),
	.w6(32'hb5596031),
	.w7(32'h36471a28),
	.w8(32'h38aece3c),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3803c9f3),
	.w1(32'h37be3322),
	.w2(32'h38a9f685),
	.w3(32'h3818abf4),
	.w4(32'h380d0d35),
	.w5(32'h38a5dd6e),
	.w6(32'h383c7f21),
	.w7(32'h385e048d),
	.w8(32'h38cc4c01),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6410028),
	.w1(32'hb73b8e9a),
	.w2(32'hb702833c),
	.w3(32'hb75a5832),
	.w4(32'hb78b4f80),
	.w5(32'hb6b50fe7),
	.w6(32'hb64f4582),
	.w7(32'hb6cb4d2e),
	.w8(32'hb5deab01),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h34e8ed81),
	.w1(32'h3500de15),
	.w2(32'hb610a0bf),
	.w3(32'h368cac8b),
	.w4(32'h360855f2),
	.w5(32'hb60363f6),
	.w6(32'h33d6017a),
	.w7(32'hb580e294),
	.w8(32'hb6897274),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5828a7e),
	.w1(32'hb797a058),
	.w2(32'hb759ffaf),
	.w3(32'h37229a12),
	.w4(32'hb78f6675),
	.w5(32'hb7144804),
	.w6(32'h36a3b21a),
	.w7(32'hb789e58d),
	.w8(32'hb6ee1152),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36cb69b0),
	.w1(32'h3776bc45),
	.w2(32'hb6cb9116),
	.w3(32'h378e47e3),
	.w4(32'h373227d7),
	.w5(32'hb767a9c7),
	.w6(32'h37c48101),
	.w7(32'h3505b051),
	.w8(32'hb7468cc2),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb86ee3d1),
	.w1(32'hb8ad2557),
	.w2(32'hb75b04cd),
	.w3(32'hb8deeab6),
	.w4(32'hb8e2a349),
	.w5(32'hb735adc9),
	.w6(32'hb7fc9d57),
	.w7(32'hb80e2058),
	.w8(32'h38246f6a),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb64b5e70),
	.w1(32'hb4682fbb),
	.w2(32'hb643163e),
	.w3(32'hb654d4b4),
	.w4(32'hb58367c1),
	.w5(32'hb698c66b),
	.w6(32'hb52da685),
	.w7(32'hb569b3cb),
	.w8(32'hb62f407f),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3732d162),
	.w1(32'h36cac4a3),
	.w2(32'hb689b7b7),
	.w3(32'h362b71c4),
	.w4(32'hb70464c1),
	.w5(32'hb7567ada),
	.w6(32'h3736e9e9),
	.w7(32'hb5deea2b),
	.w8(32'hb6878364),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb747114e),
	.w1(32'hb7797757),
	.w2(32'hb4ee6b0c),
	.w3(32'hb54f7949),
	.w4(32'hb70919ce),
	.w5(32'h377e3341),
	.w6(32'hb714a05e),
	.w7(32'hb76a79a4),
	.w8(32'h3748b935),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6e9dc95),
	.w1(32'hb6baa56f),
	.w2(32'h373cac7f),
	.w3(32'h366eaa7f),
	.w4(32'hb5827976),
	.w5(32'h37808a0a),
	.w6(32'h371d2e40),
	.w7(32'h36f73814),
	.w8(32'h37a02e43),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36e14b82),
	.w1(32'h36a2769e),
	.w2(32'h36209d51),
	.w3(32'h35147209),
	.w4(32'h35979ce6),
	.w5(32'h35af3ef1),
	.w6(32'h36d68f3c),
	.w7(32'h36210b4d),
	.w8(32'h34e1cda3),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36a13c65),
	.w1(32'h37144cb3),
	.w2(32'h370328b6),
	.w3(32'h36be6546),
	.w4(32'h36d10704),
	.w5(32'h34ae492f),
	.w6(32'h34719946),
	.w7(32'h36745ce9),
	.w8(32'hb38f3c1a),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb694d1e4),
	.w1(32'h35e3fcef),
	.w2(32'h35c5cc9a),
	.w3(32'hb69a8c4e),
	.w4(32'hb7deb415),
	.w5(32'hb7262a14),
	.w6(32'h371cc557),
	.w7(32'hb6ec8401),
	.w8(32'h37af07a3),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6d7a045),
	.w1(32'hb8b230dc),
	.w2(32'hb7ddce53),
	.w3(32'hb80c0275),
	.w4(32'hb8f50199),
	.w5(32'hb8cfec5d),
	.w6(32'h38a998c5),
	.w7(32'hb6c2fdb1),
	.w8(32'h375f999d),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38351f9c),
	.w1(32'hb70e41d7),
	.w2(32'hb7a5fda5),
	.w3(32'h3808ad9f),
	.w4(32'hb70a6ab7),
	.w5(32'hb70ccc2b),
	.w6(32'h38ecf405),
	.w7(32'h38724903),
	.w8(32'h38711dfb),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb62577e0),
	.w1(32'hb6e78397),
	.w2(32'h3514c317),
	.w3(32'hb71306a5),
	.w4(32'hb715e8c3),
	.w5(32'hb53e3a4d),
	.w6(32'hb37cf804),
	.w7(32'h357a011d),
	.w8(32'h36c36816),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h376bff47),
	.w1(32'h371e4e54),
	.w2(32'h373857b0),
	.w3(32'h3712b480),
	.w4(32'h3726932f),
	.w5(32'h369fcc94),
	.w6(32'h36764d7c),
	.w7(32'h357ed768),
	.w8(32'hb5d686b5),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb72d5446),
	.w1(32'hb5b61c45),
	.w2(32'h362e5166),
	.w3(32'hb70ac34b),
	.w4(32'h366af410),
	.w5(32'h368070de),
	.w6(32'hb62174e9),
	.w7(32'h35ff77b0),
	.w8(32'h35ad458f),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5baed8f),
	.w1(32'hb7de8098),
	.w2(32'hb7bb94a8),
	.w3(32'hb67273ab),
	.w4(32'hb8176e77),
	.w5(32'hb81c9aa3),
	.w6(32'h3723107a),
	.w7(32'hb808a369),
	.w8(32'hb7605ef3),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb81ff2bd),
	.w1(32'hb882fae0),
	.w2(32'h379ba145),
	.w3(32'hb84d9311),
	.w4(32'hb65d7119),
	.w5(32'h38839bd7),
	.w6(32'hb77eaa26),
	.w7(32'h37fc4585),
	.w8(32'h38e74181),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8691de0),
	.w1(32'hb8c699dd),
	.w2(32'hb75d5e2b),
	.w3(32'hb8a25296),
	.w4(32'hb8d50bbb),
	.w5(32'h36417a83),
	.w6(32'hb791c23c),
	.w7(32'hb7da89f9),
	.w8(32'h388cb657),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8846816),
	.w1(32'hb8bb68ee),
	.w2(32'h36ca9df0),
	.w3(32'hb8b7f919),
	.w4(32'hb8a52e9a),
	.w5(32'h381c185d),
	.w6(32'hb79341d5),
	.w7(32'hb71259d4),
	.w8(32'h38c9f70c),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb842b656),
	.w1(32'hb8695e8f),
	.w2(32'hb7ce27f2),
	.w3(32'hb888a019),
	.w4(32'hb881fdcb),
	.w5(32'h3710d4aa),
	.w6(32'h3606163e),
	.w7(32'h369489b7),
	.w8(32'h38a02f43),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb69a5e4f),
	.w1(32'h380b21f1),
	.w2(32'h38f5de7c),
	.w3(32'h36fe2d07),
	.w4(32'h38056f6c),
	.w5(32'h38ca3d90),
	.w6(32'hb6451347),
	.w7(32'h382c60eb),
	.w8(32'h38d389a9),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36a3822a),
	.w1(32'h35c3acab),
	.w2(32'hb71f631a),
	.w3(32'hb7411f0a),
	.w4(32'hb6fe742e),
	.w5(32'hb692864d),
	.w6(32'hb7003abb),
	.w7(32'h34147fe7),
	.w8(32'h372640e2),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb82625ac),
	.w1(32'hb74f3551),
	.w2(32'h37ecb1b3),
	.w3(32'hb8305fa1),
	.w4(32'hb7466c22),
	.w5(32'h37ceb445),
	.w6(32'hb6f88996),
	.w7(32'h37bcc56d),
	.w8(32'h38613fda),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb78acb3b),
	.w1(32'h37694257),
	.w2(32'h3828e3a7),
	.w3(32'hb7ea6b25),
	.w4(32'h368801f1),
	.w5(32'h3807d784),
	.w6(32'hb7d318c1),
	.w7(32'h3724b26b),
	.w8(32'h37de4b68),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h371bea1b),
	.w1(32'hb7a9b140),
	.w2(32'h37343f93),
	.w3(32'hb53638a2),
	.w4(32'hb70f2bb4),
	.w5(32'h377f6d40),
	.w6(32'h356238d9),
	.w7(32'hb72f56da),
	.w8(32'h3733575b),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb270927b),
	.w1(32'h368caf2d),
	.w2(32'h373df10d),
	.w3(32'h364ab10a),
	.w4(32'h36d70269),
	.w5(32'h373f67f8),
	.w6(32'h36b3707e),
	.w7(32'h36ea5177),
	.w8(32'h37413a62),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb71fb0d8),
	.w1(32'hb7a54a71),
	.w2(32'h37c68a7b),
	.w3(32'h36d11040),
	.w4(32'h378acb79),
	.w5(32'h38795813),
	.w6(32'hb6d66780),
	.w7(32'h35207bdb),
	.w8(32'h380de26b),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h374b32bd),
	.w1(32'h372e9dde),
	.w2(32'h36df0505),
	.w3(32'h3748a418),
	.w4(32'h36ee57c3),
	.w5(32'h364e906f),
	.w6(32'h37496af2),
	.w7(32'h36dc08b4),
	.w8(32'h3668db6c),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5f89806),
	.w1(32'hb4b95574),
	.w2(32'h34d2599d),
	.w3(32'hb57a7d7b),
	.w4(32'h34bb6138),
	.w5(32'h35c2e0db),
	.w6(32'h3499f5d6),
	.w7(32'hb524e4ad),
	.w8(32'hb514a7c4),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb60d250f),
	.w1(32'h34e242cd),
	.w2(32'h349a0771),
	.w3(32'hb6037bba),
	.w4(32'h35b2fc84),
	.w5(32'h35ac0d24),
	.w6(32'hb4cef4f1),
	.w7(32'hb4b2787f),
	.w8(32'hb591a9a5),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb53538c9),
	.w1(32'hb5ee8eca),
	.w2(32'hb55e4e81),
	.w3(32'hb564abf7),
	.w4(32'hb622bc90),
	.w5(32'hb68618a5),
	.w6(32'hb5e88ba7),
	.w7(32'hb5614921),
	.w8(32'hb62cc6f9),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb74adc4d),
	.w1(32'hb7bb5a72),
	.w2(32'hb7663a7e),
	.w3(32'hb74aaff4),
	.w4(32'hb791f525),
	.w5(32'hb7717113),
	.w6(32'h3725459e),
	.w7(32'hb5508194),
	.w8(32'h37827870),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h364996ad),
	.w1(32'hb75dcd62),
	.w2(32'hb7577c01),
	.w3(32'hb66bd473),
	.w4(32'hb6b67fb1),
	.w5(32'hb6a81578),
	.w6(32'h35c4234a),
	.w7(32'h3694916c),
	.w8(32'h36e42f26),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h371267e6),
	.w1(32'h363b2d09),
	.w2(32'h37c62449),
	.w3(32'h37283358),
	.w4(32'h3735acc3),
	.w5(32'h37c6f3cf),
	.w6(32'h3729e2d3),
	.w7(32'h374e64bb),
	.w8(32'h37ae129d),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h379368b0),
	.w1(32'hb6901ca6),
	.w2(32'hb68c57ad),
	.w3(32'h37eef902),
	.w4(32'hb5a91cd3),
	.w5(32'hb6049e07),
	.w6(32'h37a8277f),
	.w7(32'hb6486e0b),
	.w8(32'hb6357978),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb604e20c),
	.w1(32'hb5c7016c),
	.w2(32'h35e16f49),
	.w3(32'hb6a34c6c),
	.w4(32'hb6defc78),
	.w5(32'hb5ce5ff1),
	.w6(32'hb614c151),
	.w7(32'hb684547a),
	.w8(32'hb5dcfd58),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb48659ff),
	.w1(32'h34f238e8),
	.w2(32'hb475aff5),
	.w3(32'h354bfac5),
	.w4(32'h3520754d),
	.w5(32'h34c504d6),
	.w6(32'hb580d7f5),
	.w7(32'hb58974e0),
	.w8(32'hb5edd447),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5f59558),
	.w1(32'hb6640bcb),
	.w2(32'hb6f6d6f4),
	.w3(32'h36700b92),
	.w4(32'hb660de47),
	.w5(32'hb6ba84d8),
	.w6(32'h340af602),
	.w7(32'hb65839ca),
	.w8(32'hb5c33a8b),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35895d3c),
	.w1(32'h34f6cde4),
	.w2(32'hb5a1b03e),
	.w3(32'h35c3bfcf),
	.w4(32'hb4c012e4),
	.w5(32'hb6189dae),
	.w6(32'h34980e72),
	.w7(32'hb5941764),
	.w8(32'hb6771503),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37db4624),
	.w1(32'h37292b70),
	.w2(32'hb72b8325),
	.w3(32'h37b7f7f1),
	.w4(32'h37f79f11),
	.w5(32'h379dad45),
	.w6(32'h37d651b6),
	.w7(32'h3562a626),
	.w8(32'hb75158f3),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37af3a3f),
	.w1(32'h36e7aa65),
	.w2(32'h381d5bb7),
	.w3(32'h3762366c),
	.w4(32'h3737784f),
	.w5(32'h38635827),
	.w6(32'h3838bb8b),
	.w7(32'h382e5fff),
	.w8(32'h38ad3ab2),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37e7963f),
	.w1(32'h372455e0),
	.w2(32'h37e0ffa6),
	.w3(32'h381b2596),
	.w4(32'h373085ea),
	.w5(32'h37acb0cc),
	.w6(32'h3898ef91),
	.w7(32'h38305722),
	.w8(32'h3871861b),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3736792f),
	.w1(32'hb7f224a6),
	.w2(32'h386f2384),
	.w3(32'hb811db29),
	.w4(32'hb88719a1),
	.w5(32'h37f281ca),
	.w6(32'h3808a982),
	.w7(32'hb4e92c10),
	.w8(32'h38dbd734),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h350e79de),
	.w1(32'h33bf981f),
	.w2(32'hb598e383),
	.w3(32'hb5283ca5),
	.w4(32'h31750e34),
	.w5(32'hb5a846e5),
	.w6(32'hb5e48b37),
	.w7(32'hb5a81db5),
	.w8(32'hb627c9ad),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb4b516ee),
	.w1(32'hb4b1b59f),
	.w2(32'hb60a223c),
	.w3(32'hb49e5c53),
	.w4(32'hb4e78340),
	.w5(32'hb6158404),
	.w6(32'hb6747965),
	.w7(32'hb628bd8a),
	.w8(32'hb6913cc5),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5735382),
	.w1(32'hb5ebd78b),
	.w2(32'hb64dc183),
	.w3(32'hb60e7464),
	.w4(32'hb54d08fc),
	.w5(32'hb5c4b1b1),
	.w6(32'hb68091ac),
	.w7(32'hb61bf71b),
	.w8(32'hb625d2bc),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3770107a),
	.w1(32'h371f387a),
	.w2(32'h36e64a11),
	.w3(32'h378c44b0),
	.w4(32'h37146d34),
	.w5(32'h373c92ba),
	.w6(32'h3736f671),
	.w7(32'h37312ce7),
	.w8(32'h36a0c7f7),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6be059d),
	.w1(32'h34ef609c),
	.w2(32'h364d2b2a),
	.w3(32'hb7063c51),
	.w4(32'hb6941bcd),
	.w5(32'hb4facd6f),
	.w6(32'hb6ec5c1a),
	.w7(32'hb5acab03),
	.w8(32'h3686a67b),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36cfb630),
	.w1(32'h37334ef6),
	.w2(32'h3788ff63),
	.w3(32'h375dbf14),
	.w4(32'h37beac5c),
	.w5(32'h37b69fa6),
	.w6(32'h3683654d),
	.w7(32'h36c3267e),
	.w8(32'h35e1921c),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h379bbd59),
	.w1(32'h3819c2ed),
	.w2(32'h385830c3),
	.w3(32'hb4b756db),
	.w4(32'h37eb9b2b),
	.w5(32'h38331a7a),
	.w6(32'h378ac789),
	.w7(32'h3820f840),
	.w8(32'h38327c9a),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7d1984d),
	.w1(32'hb7cac737),
	.w2(32'h3841b816),
	.w3(32'hb8321abd),
	.w4(32'hb7f8a35c),
	.w5(32'h383b674a),
	.w6(32'hb7db5d46),
	.w7(32'hb70801f5),
	.w8(32'h386f2e25),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37501049),
	.w1(32'hb68700d4),
	.w2(32'h37c00527),
	.w3(32'h3719d07a),
	.w4(32'hb5961932),
	.w5(32'h37cd4ed9),
	.w6(32'h378b45e5),
	.w7(32'h369b37dc),
	.w8(32'h38033014),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35d6ba8f),
	.w1(32'hb6e30558),
	.w2(32'h37061d98),
	.w3(32'h3688b011),
	.w4(32'h37230e5c),
	.w5(32'h380b82ae),
	.w6(32'h369fefcb),
	.w7(32'hb57047e1),
	.w8(32'h3780ca9a),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6deee7a),
	.w1(32'hb75dda76),
	.w2(32'h3720931b),
	.w3(32'hb6453313),
	.w4(32'hb68f8635),
	.w5(32'h377657e9),
	.w6(32'h3735f9e2),
	.w7(32'h3678a352),
	.w8(32'h37aa1fd6),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb623219a),
	.w1(32'hb60f8955),
	.w2(32'h37a558f2),
	.w3(32'h3609b6b9),
	.w4(32'h373cee60),
	.w5(32'h3819fd89),
	.w6(32'h367a6363),
	.w7(32'h37395a83),
	.w8(32'h38080b51),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h34aebc2c),
	.w1(32'h34f2398a),
	.w2(32'hb4512b46),
	.w3(32'h3514da87),
	.w4(32'h33ddac24),
	.w5(32'h33e6b929),
	.w6(32'h34b81af1),
	.w7(32'h3396e15a),
	.w8(32'hb4126c2f),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb53e458d),
	.w1(32'hb55fe771),
	.w2(32'hb5b6e572),
	.w3(32'hb54264cf),
	.w4(32'hb51b3819),
	.w5(32'hb588643e),
	.w6(32'hb5a48e1a),
	.w7(32'hb545273e),
	.w8(32'hb4111eda),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb395cbbc),
	.w1(32'h330d9854),
	.w2(32'h361e5509),
	.w3(32'hb360f0a9),
	.w4(32'hb42bb6ab),
	.w5(32'h35573c82),
	.w6(32'hb4e4135b),
	.w7(32'h3325e7e9),
	.w8(32'hb653c084),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5fc9856),
	.w1(32'hb5337056),
	.w2(32'h358dcec9),
	.w3(32'hb65832d3),
	.w4(32'hb54c39da),
	.w5(32'h34a9f9b6),
	.w6(32'hb50d0d38),
	.w7(32'hb54014f7),
	.w8(32'hb44d99fc),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37f1fa32),
	.w1(32'hb6dcf28c),
	.w2(32'hb796a6a0),
	.w3(32'h37c928ee),
	.w4(32'hb65eebac),
	.w5(32'hb718ed9e),
	.w6(32'h37ae1010),
	.w7(32'hb73cdac9),
	.w8(32'h340d90ee),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h360d249d),
	.w1(32'h3611b818),
	.w2(32'hb5e02b69),
	.w3(32'hb603e249),
	.w4(32'hb69afb01),
	.w5(32'hb6ca4b85),
	.w6(32'h37050b0c),
	.w7(32'h36851bd6),
	.w8(32'h36207c9a),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb787cc0b),
	.w1(32'hb7f65f99),
	.w2(32'h378d560a),
	.w3(32'hb7ee816d),
	.w4(32'hb76e79b9),
	.w5(32'h380faedd),
	.w6(32'hb789d6b2),
	.w7(32'h354721da),
	.w8(32'h3834034f),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37f14134),
	.w1(32'h377b6c5f),
	.w2(32'h3808e61a),
	.w3(32'h3845f894),
	.w4(32'h37ad7e37),
	.w5(32'h38287b3b),
	.w6(32'h381ac996),
	.w7(32'h381f1016),
	.w8(32'h38355a07),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37ce8a38),
	.w1(32'hb75449a4),
	.w2(32'hb755ceee),
	.w3(32'h37abcc4f),
	.w4(32'hb7c3fab0),
	.w5(32'hb7ef604f),
	.w6(32'h381dd3f1),
	.w7(32'hb74f8bd1),
	.w8(32'hb64dd001),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38372250),
	.w1(32'hb6e0a377),
	.w2(32'h37a9f802),
	.w3(32'h3828da11),
	.w4(32'h37e1b52c),
	.w5(32'h3831931f),
	.w6(32'h37e8f7bd),
	.w7(32'h376a67cc),
	.w8(32'h38079b60),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7d28761),
	.w1(32'hb820741a),
	.w2(32'hb7547810),
	.w3(32'hb7c337c1),
	.w4(32'hb81d4626),
	.w5(32'hb74a2564),
	.w6(32'h378aa83c),
	.w7(32'hb6d59032),
	.w8(32'h37b8fcd2),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h379c7190),
	.w1(32'hb7748b93),
	.w2(32'h37907062),
	.w3(32'h370ee502),
	.w4(32'hb7c78ea1),
	.w5(32'h37acfbee),
	.w6(32'h379633bf),
	.w7(32'hb72e3df3),
	.w8(32'h37f16a6c),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb76d1bf0),
	.w1(32'hb7cabd74),
	.w2(32'hb72074a9),
	.w3(32'hb7435083),
	.w4(32'hb576173f),
	.w5(32'h3785a38b),
	.w6(32'h36b1d4f6),
	.w7(32'hb5179a63),
	.w8(32'h379703ca),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6895533),
	.w1(32'hb7d69e84),
	.w2(32'h37625323),
	.w3(32'hb74a6409),
	.w4(32'hb81533ad),
	.w5(32'h36c16261),
	.w6(32'h36c71adf),
	.w7(32'hb788ef96),
	.w8(32'h378b978f),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb81a7062),
	.w1(32'hb820993f),
	.w2(32'h368aca0f),
	.w3(32'hb6ea3d4e),
	.w4(32'hb6db6e33),
	.w5(32'h37983fdd),
	.w6(32'hb7963005),
	.w7(32'hb713fb2e),
	.w8(32'h3743c221),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f69324),
	.w1(32'hb8ffb79d),
	.w2(32'h3813bd49),
	.w3(32'hb87af47b),
	.w4(32'hb7e8df1c),
	.w5(32'h38833027),
	.w6(32'hb7b5508c),
	.w7(32'h3773a7dd),
	.w8(32'h38cfa3a9),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb85d66d0),
	.w1(32'hb848226c),
	.w2(32'hb7e2bd8b),
	.w3(32'hb83406d6),
	.w4(32'hb813a6a6),
	.w5(32'h3771fbb6),
	.w6(32'h385aecbe),
	.w7(32'h389d3198),
	.w8(32'h38f716c0),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37b63895),
	.w1(32'h3868e784),
	.w2(32'h38bf0285),
	.w3(32'h382738f2),
	.w4(32'h38a1864e),
	.w5(32'h388f54f2),
	.w6(32'h3790ce68),
	.w7(32'h38564b0e),
	.w8(32'h387ff21b),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38050818),
	.w1(32'hb912bb1a),
	.w2(32'hb8b588e4),
	.w3(32'hb8972aa7),
	.w4(32'hb91c59bc),
	.w5(32'hb89df974),
	.w6(32'h389b028f),
	.w7(32'hb75c6229),
	.w8(32'h38b68904),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89d9fe5),
	.w1(32'hb8a359ff),
	.w2(32'h38695e53),
	.w3(32'hb891875f),
	.w4(32'hb81abb50),
	.w5(32'h3887159e),
	.w6(32'hb7627a13),
	.w7(32'h361db4e1),
	.w8(32'h38de87ce),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6df3b95),
	.w1(32'hb7ce8beb),
	.w2(32'h34e0e1c0),
	.w3(32'hb79f6636),
	.w4(32'hb783f625),
	.w5(32'h375dcb69),
	.w6(32'hb706fc9f),
	.w7(32'hb722d07f),
	.w8(32'h37c83b3f),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7ac7b3a),
	.w1(32'hb7ca51e9),
	.w2(32'h38232d31),
	.w3(32'hb8ba2097),
	.w4(32'hb7f6c583),
	.w5(32'h370d058f),
	.w6(32'hb7dec748),
	.w7(32'hb69156c3),
	.w8(32'h3864e7e0),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37a4c173),
	.w1(32'h37f8afa1),
	.w2(32'h3891aa39),
	.w3(32'h3795b61f),
	.w4(32'h382f2002),
	.w5(32'h38b7dc64),
	.w6(32'h35396eec),
	.w7(32'h37bf88a1),
	.w8(32'h37f0f5ad),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35ec2141),
	.w1(32'hb6ba7f93),
	.w2(32'hb7cd0ba0),
	.w3(32'hb6bfc45f),
	.w4(32'hb72f405f),
	.w5(32'hb779337c),
	.w6(32'hb3fe80b5),
	.w7(32'hb707f2ad),
	.w8(32'hb6282438),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35ef17e3),
	.w1(32'h3592256e),
	.w2(32'h35533c5e),
	.w3(32'h35e08b00),
	.w4(32'h369584aa),
	.w5(32'h369e112d),
	.w6(32'h36da0c8f),
	.w7(32'h3705c0a1),
	.w8(32'h370c3eae),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36000f35),
	.w1(32'hb725144d),
	.w2(32'hb64ba07f),
	.w3(32'hb781fb82),
	.w4(32'hb74e1b86),
	.w5(32'hb70c6759),
	.w6(32'hb66ce8a3),
	.w7(32'hb63164de),
	.w8(32'h36372988),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb85da202),
	.w1(32'hb7d458a6),
	.w2(32'h38136613),
	.w3(32'hb7d00fd1),
	.w4(32'h37c6570a),
	.w5(32'h38c399b4),
	.w6(32'hb7acc7ba),
	.w7(32'h3792bfc7),
	.w8(32'h38a3e5d4),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88f0291),
	.w1(32'hb8c84e8c),
	.w2(32'h35ddcfd1),
	.w3(32'hb886ceed),
	.w4(32'hb848c54a),
	.w5(32'h3766cdda),
	.w6(32'hb7df4e23),
	.w7(32'hb801575c),
	.w8(32'h384e4e40),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36e53a80),
	.w1(32'hb7da256e),
	.w2(32'hb67d6bbe),
	.w3(32'hb7a1fa17),
	.w4(32'hb83a94e9),
	.w5(32'hb79b2116),
	.w6(32'h37301153),
	.w7(32'hb7a5c248),
	.w8(32'h360febb5),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb77e524f),
	.w1(32'hb81613ff),
	.w2(32'hb6b731a4),
	.w3(32'hb8295fe2),
	.w4(32'hb809b3f9),
	.w5(32'h34d5532c),
	.w6(32'hb7049dcd),
	.w7(32'hb74c64c2),
	.w8(32'h37d35ff2),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3809bcc4),
	.w1(32'h37cb7c2a),
	.w2(32'h3786ec3d),
	.w3(32'h3765a02a),
	.w4(32'hb5fd710f),
	.w5(32'hb68f19d3),
	.w6(32'h376baf39),
	.w7(32'h35d94ace),
	.w8(32'h3717aa83),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7ba0532),
	.w1(32'hb815ce05),
	.w2(32'h368cb236),
	.w3(32'hb76ec5ac),
	.w4(32'hb7c71b37),
	.w5(32'h3643a996),
	.w6(32'h379e5ba8),
	.w7(32'h36a5ad9c),
	.w8(32'h37f8c7c0),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7543d02),
	.w1(32'hb7d83c8e),
	.w2(32'h36b39415),
	.w3(32'hb71d8d0a),
	.w4(32'hb71b52d8),
	.w5(32'h37d04c8e),
	.w6(32'h35fd4329),
	.w7(32'h36ccb0d6),
	.w8(32'h381e1df3),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h35866cf2),
	.w1(32'h35b44936),
	.w2(32'h3564a3d0),
	.w3(32'h35cb17e3),
	.w4(32'h350bec10),
	.w5(32'h364e434e),
	.w6(32'hb629edbe),
	.w7(32'hb5796995),
	.w8(32'h344aa0af),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h341c0d80),
	.w1(32'hb4617ee6),
	.w2(32'hb59c2c70),
	.w3(32'hb48439fa),
	.w4(32'h3573d907),
	.w5(32'h34bb6e6e),
	.w6(32'hb4fc44cb),
	.w7(32'hb4f6211e),
	.w8(32'hb5af3c5c),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb59c2058),
	.w1(32'hb58ab00f),
	.w2(32'hb53d87b9),
	.w3(32'hb5067bbc),
	.w4(32'hb5223795),
	.w5(32'hb5c3c59f),
	.w6(32'hb5526d17),
	.w7(32'hb51909c3),
	.w8(32'hb595bda9),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3686afce),
	.w1(32'h36a2f928),
	.w2(32'h36c9aaec),
	.w3(32'h3626fe90),
	.w4(32'h35c3efe7),
	.w5(32'h36b520fd),
	.w6(32'h354ae3d8),
	.w7(32'hb58191c1),
	.w8(32'h3514bcbe),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb80aa472),
	.w1(32'hb852c198),
	.w2(32'h36a1e022),
	.w3(32'hb810c3dc),
	.w4(32'hb81005e0),
	.w5(32'h37ad3112),
	.w6(32'hb754d977),
	.w7(32'hb742b983),
	.w8(32'h37ff2ecb),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3726feb4),
	.w1(32'hb65ffa95),
	.w2(32'hb63a4d72),
	.w3(32'h365cc3d5),
	.w4(32'hb6fe20fd),
	.w5(32'h35c3a1ce),
	.w6(32'h3493cd7f),
	.w7(32'hb70031eb),
	.w8(32'hb4d41ba7),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h362c5a63),
	.w1(32'h3662232d),
	.w2(32'h374822b3),
	.w3(32'hb509b9da),
	.w4(32'h36d26d16),
	.w5(32'h3783e302),
	.w6(32'hb608cea0),
	.w7(32'h366aed84),
	.w8(32'h37395444),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h379d76be),
	.w1(32'h35b98fe1),
	.w2(32'h3796b928),
	.w3(32'h36e518ab),
	.w4(32'hb581022f),
	.w5(32'h379f2fb5),
	.w6(32'h37952528),
	.w7(32'h3742a9d7),
	.w8(32'h381c0547),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb4d8e630),
	.w1(32'hb578ea64),
	.w2(32'hb60fe42d),
	.w3(32'hb5742bdd),
	.w4(32'h356afe29),
	.w5(32'hb541ef8e),
	.w6(32'hb5aabf7d),
	.w7(32'hb582016f),
	.w8(32'hb5e343a2),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h365f97fe),
	.w1(32'h3638eb38),
	.w2(32'h369a2036),
	.w3(32'hb4c481e1),
	.w4(32'h35ee591a),
	.w5(32'h3608454e),
	.w6(32'h3685fc7d),
	.w7(32'h365d20cd),
	.w8(32'h366dc129),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h332ccef7),
	.w1(32'h353722f9),
	.w2(32'hb56bf3ab),
	.w3(32'hb68f7840),
	.w4(32'hb61a99ac),
	.w5(32'hb68e3263),
	.w6(32'hb48fdc29),
	.w7(32'hb5081426),
	.w8(32'hb51b8648),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb701cf6a),
	.w1(32'hbbb6e7ed),
	.w2(32'hba73d06e),
	.w3(32'hb76e5135),
	.w4(32'hbc3700ae),
	.w5(32'hbc2a753a),
	.w6(32'hb9b1b54d),
	.w7(32'h3c2f88a6),
	.w8(32'hba1c9541),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4ff9a9),
	.w1(32'hbb15e8ab),
	.w2(32'h3b861e75),
	.w3(32'hbbc14ac1),
	.w4(32'hbb5608ba),
	.w5(32'hbb0d02dd),
	.w6(32'h39d244de),
	.w7(32'h3c301523),
	.w8(32'hbaac4c4e),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8da9b03),
	.w1(32'hbc70efdc),
	.w2(32'hbc750c26),
	.w3(32'h39e99cf2),
	.w4(32'h3bc86e12),
	.w5(32'h3b770063),
	.w6(32'hbc7ca0fb),
	.w7(32'hbbcbd227),
	.w8(32'h3b28e47a),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc150500),
	.w1(32'hb92aa2f7),
	.w2(32'h3bb1d551),
	.w3(32'hbbe98453),
	.w4(32'h3c41b84e),
	.w5(32'h3cd6aead),
	.w6(32'hbc238242),
	.w7(32'hbc922d2a),
	.w8(32'hbbed1e12),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baa93df),
	.w1(32'hbbc586a5),
	.w2(32'hba1ac394),
	.w3(32'h3c4c5d57),
	.w4(32'h3a9cdbdb),
	.w5(32'h3be0e659),
	.w6(32'hbbd7da6b),
	.w7(32'hbc093007),
	.w8(32'hba756adf),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb455bae),
	.w1(32'hbc3e80ad),
	.w2(32'hbb2e160d),
	.w3(32'h3b8ea030),
	.w4(32'hba16f450),
	.w5(32'h3c899a28),
	.w6(32'hbc0fa646),
	.w7(32'hbc0b0ed7),
	.w8(32'hbc1cbd9d),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc314c68),
	.w1(32'h3ba27e7f),
	.w2(32'hbbf739fc),
	.w3(32'h3b197f19),
	.w4(32'hbb955a0d),
	.w5(32'hbc0ed694),
	.w6(32'h3c3e4f33),
	.w7(32'hbb483bcd),
	.w8(32'hbc0743f2),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc07721),
	.w1(32'hbb0109ed),
	.w2(32'h39ade388),
	.w3(32'h3c22ec9f),
	.w4(32'h3abfa6d3),
	.w5(32'h3bbec6b6),
	.w6(32'hbab500b1),
	.w7(32'h3bacb20b),
	.w8(32'hbb2d31dd),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeb5dec),
	.w1(32'hbbea34bc),
	.w2(32'hb7c4067e),
	.w3(32'h3c463d13),
	.w4(32'h3b924734),
	.w5(32'h3c87bdb6),
	.w6(32'hbc67da3b),
	.w7(32'hbcc71023),
	.w8(32'hbc378403),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab43040),
	.w1(32'h398af2a4),
	.w2(32'h3bc3e7b1),
	.w3(32'h3c100f94),
	.w4(32'hbbec802f),
	.w5(32'hbc2dfe8d),
	.w6(32'h3bb27103),
	.w7(32'h3ca66bc8),
	.w8(32'h3b4e57fa),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba00a88d),
	.w1(32'hbb2f8598),
	.w2(32'h3a987984),
	.w3(32'hbbb0cc90),
	.w4(32'hbbb99f8b),
	.w5(32'hbb807778),
	.w6(32'hbb558a52),
	.w7(32'h3b855db8),
	.w8(32'hba9907de),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab96e2a),
	.w1(32'hbbc4d533),
	.w2(32'hbbfd43d6),
	.w3(32'h386b5cb1),
	.w4(32'h3c8dabf6),
	.w5(32'h3d11d703),
	.w6(32'hbc776a31),
	.w7(32'hbd057bf7),
	.w8(32'hbc2bd06e),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb906b612),
	.w1(32'hbcadc264),
	.w2(32'hbcb9bf61),
	.w3(32'h3c93bc57),
	.w4(32'hba950213),
	.w5(32'h3b68052e),
	.w6(32'hbb7f4544),
	.w7(32'hbb28f315),
	.w8(32'hbbcc9454),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb37701),
	.w1(32'h3b8ff097),
	.w2(32'h3c6bbc75),
	.w3(32'hb7f6a6f9),
	.w4(32'h3b0e1427),
	.w5(32'h3b838736),
	.w6(32'h3b978ceb),
	.w7(32'h3c1bee71),
	.w8(32'h3bfbd2ba),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bec77a1),
	.w1(32'hbb494b82),
	.w2(32'hbb256422),
	.w3(32'h3bfa2ef3),
	.w4(32'hbbe28a69),
	.w5(32'hbc068b7a),
	.w6(32'hbb26067d),
	.w7(32'h3b93ae1c),
	.w8(32'hbaa911d7),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7db1e7),
	.w1(32'hba957c67),
	.w2(32'h3bbce80c),
	.w3(32'hbba0869e),
	.w4(32'hbc60edc1),
	.w5(32'hbcc8ceee),
	.w6(32'h3c2c93b5),
	.w7(32'h3cee4546),
	.w8(32'h3b3ff25d),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b4594),
	.w1(32'h3bbe7e9c),
	.w2(32'h3c47cf2c),
	.w3(32'hbc9fbb31),
	.w4(32'hba7f40bf),
	.w5(32'h3ab2125e),
	.w6(32'h3b299e83),
	.w7(32'hbb9a1012),
	.w8(32'h3aa6df2d),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1de355),
	.w1(32'h397cd4d9),
	.w2(32'h3b369723),
	.w3(32'h3b0fbfbe),
	.w4(32'hba66d7db),
	.w5(32'h3890dd2b),
	.w6(32'hbb3aa281),
	.w7(32'h3b078c10),
	.w8(32'hba8502c9),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1ca934),
	.w1(32'hbaf7ec80),
	.w2(32'h3b0c7e60),
	.w3(32'hb7da72d5),
	.w4(32'hbba02bfc),
	.w5(32'hbc231547),
	.w6(32'hbb873bf3),
	.w7(32'h3a2f4bbf),
	.w8(32'h391fd6d1),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b365626),
	.w1(32'hbbf46a18),
	.w2(32'hbb7b67b8),
	.w3(32'h3a03f908),
	.w4(32'h3c32c50e),
	.w5(32'h3ce70f0c),
	.w6(32'hbca0f179),
	.w7(32'hbd0ebc4b),
	.w8(32'hbc6403bb),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39868f47),
	.w1(32'hb90b5803),
	.w2(32'h3bc45a56),
	.w3(32'h3c4040a6),
	.w4(32'h3b951e39),
	.w5(32'h3c716fe2),
	.w6(32'hbbf10a63),
	.w7(32'hbc289b60),
	.w8(32'hbb7651fa),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5c358e),
	.w1(32'hbae3f4ec),
	.w2(32'hb8f5c9ca),
	.w3(32'h3bb66522),
	.w4(32'hbb595eb3),
	.w5(32'hbb077aeb),
	.w6(32'hbb159da2),
	.w7(32'h3a7ca52a),
	.w8(32'hbaa7ee5a),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a74329a),
	.w1(32'hbc851f5f),
	.w2(32'hbc2b7f53),
	.w3(32'hb9937728),
	.w4(32'hbc1a2176),
	.w5(32'hbc108fce),
	.w6(32'hbbee7fe9),
	.w7(32'h3bd3b720),
	.w8(32'hbb049710),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0fcb9a),
	.w1(32'hbc970371),
	.w2(32'hbc3fe3f5),
	.w3(32'hbb9c5340),
	.w4(32'hbac9934b),
	.w5(32'hbc920a03),
	.w6(32'hbbce3a19),
	.w7(32'hbba92150),
	.w8(32'hbb7b1617),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcacd13a),
	.w1(32'hbb9e059f),
	.w2(32'hbbad530f),
	.w3(32'hbb8741b5),
	.w4(32'hbb445b5e),
	.w5(32'hbb18e55c),
	.w6(32'hbb831de6),
	.w7(32'hbab0520f),
	.w8(32'hbafee7e7),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac4d1a0),
	.w1(32'hbaa8fcbc),
	.w2(32'h3bb79282),
	.w3(32'h3b181ffa),
	.w4(32'hbbdd1a68),
	.w5(32'hbc0c6cf5),
	.w6(32'h3b889376),
	.w7(32'h3c9ae5ba),
	.w8(32'h3afdf320),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaecb934),
	.w1(32'h3b02c5c3),
	.w2(32'h3be80669),
	.w3(32'hbbaa979b),
	.w4(32'h3bb3ed6e),
	.w5(32'h3c3656ef),
	.w6(32'hbbcdd02a),
	.w7(32'hbc0e94e8),
	.w8(32'hba5c4a6b),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1babb1),
	.w1(32'hbc0dc1c6),
	.w2(32'h3a68dbdb),
	.w3(32'h3ad5f26e),
	.w4(32'hbba9cf2e),
	.w5(32'hbc45093f),
	.w6(32'h3b442a65),
	.w7(32'h3c598ba6),
	.w8(32'h3b47664d),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc17df4a),
	.w1(32'hbbb6c0f8),
	.w2(32'hbb5dc884),
	.w3(32'hbbb1f286),
	.w4(32'hbbeb3805),
	.w5(32'hbbe2cbb9),
	.w6(32'hbb830de7),
	.w7(32'h3a06eed6),
	.w8(32'hbb740f3a),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7f368c),
	.w1(32'hbbba4448),
	.w2(32'h3b524e68),
	.w3(32'hbb551237),
	.w4(32'h3c0718f3),
	.w5(32'h3c45dab8),
	.w6(32'hbc5c345a),
	.w7(32'hbc06c612),
	.w8(32'hba8b8101),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb818497),
	.w1(32'hbc24fef0),
	.w2(32'hbbea895d),
	.w3(32'hbc08ee4c),
	.w4(32'hbb801051),
	.w5(32'hba86035c),
	.w6(32'hbc230c40),
	.w7(32'hbbd22170),
	.w8(32'hbb9da9c6),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb656c9d),
	.w1(32'hbba55754),
	.w2(32'hbb547c32),
	.w3(32'h3b338a37),
	.w4(32'hbae2dfdd),
	.w5(32'hbae25494),
	.w6(32'hbbe3eb5d),
	.w7(32'hbae8dbc9),
	.w8(32'h3a5c617a),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a09184),
	.w1(32'hbbf9dd79),
	.w2(32'hbbb92f04),
	.w3(32'h3ab21697),
	.w4(32'hbbe48691),
	.w5(32'hbbd6f158),
	.w6(32'hbbb8e377),
	.w7(32'h3abef314),
	.w8(32'hbb6954b1),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba34b3a),
	.w1(32'hbc0ed801),
	.w2(32'hbbf3a3a9),
	.w3(32'hbb429f65),
	.w4(32'hbc02e67a),
	.w5(32'hbc0964f0),
	.w6(32'hbba96ef8),
	.w7(32'hb9b30e55),
	.w8(32'hbbd31c85),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbff0603),
	.w1(32'h3a4c48c2),
	.w2(32'h3a2f99a6),
	.w3(32'hbbaf45aa),
	.w4(32'h3a19fe29),
	.w5(32'hbb8b4eaa),
	.w6(32'hbb8b455e),
	.w7(32'hba892e0a),
	.w8(32'h3833e5ee),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0f9fcc),
	.w1(32'h3aa28454),
	.w2(32'h3b8c90c3),
	.w3(32'hbb8ef28e),
	.w4(32'hbc18c2ac),
	.w5(32'hbbcb0018),
	.w6(32'h3b1d7c1c),
	.w7(32'hbb724330),
	.w8(32'hbb8e42e5),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba934e2),
	.w1(32'hbc35f8e7),
	.w2(32'hbc4665c2),
	.w3(32'hbc07139d),
	.w4(32'h3c661931),
	.w5(32'h3d0cfbec),
	.w6(32'hbcb2eea8),
	.w7(32'hbd017c9f),
	.w8(32'hbc2f1de5),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b23de98),
	.w1(32'hbbe391fb),
	.w2(32'hbb8a1d41),
	.w3(32'h3c9f607d),
	.w4(32'hbba9a15f),
	.w5(32'hbaf64444),
	.w6(32'hbb9ee818),
	.w7(32'hba1f5f1a),
	.w8(32'hbb1b8c2a),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8707f3),
	.w1(32'h3acbd7e5),
	.w2(32'h3bca6022),
	.w3(32'h3a9819bb),
	.w4(32'h3c28e5f1),
	.w5(32'h3ce54163),
	.w6(32'hbc1eb6e4),
	.w7(32'hbcad5dcf),
	.w8(32'hbbf8fc10),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c18bdfb),
	.w1(32'hbb8e19dc),
	.w2(32'h3a83f964),
	.w3(32'h3c9826c3),
	.w4(32'h3bc2a8eb),
	.w5(32'h3c8e9051),
	.w6(32'hbc3d5c6d),
	.w7(32'hbca51fce),
	.w8(32'hbc100138),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395fb964),
	.w1(32'hbb9eec8d),
	.w2(32'h3b07bd45),
	.w3(32'h3c0a9730),
	.w4(32'hbbc08fad),
	.w5(32'hbbdb0ca8),
	.w6(32'hba765342),
	.w7(32'h3c479e85),
	.w8(32'hba9eb2d7),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb21a912),
	.w1(32'hbb0a19cc),
	.w2(32'h3b7e7344),
	.w3(32'hbb55723b),
	.w4(32'hb97711ad),
	.w5(32'h3c4acaef),
	.w6(32'hbc27eed3),
	.w7(32'hbc852a5e),
	.w8(32'hbbf50881),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b94fed3),
	.w1(32'hbb1cc427),
	.w2(32'hbbd260e5),
	.w3(32'h3bc79c03),
	.w4(32'hbad5a2ae),
	.w5(32'hbb986b57),
	.w6(32'hbb48cf08),
	.w7(32'hbb0ede94),
	.w8(32'h3b135151),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a216b9),
	.w1(32'hbaad5cc7),
	.w2(32'h3ba8ce9b),
	.w3(32'h3a680b91),
	.w4(32'hbae6ea4d),
	.w5(32'h3c262260),
	.w6(32'hbbcfbff0),
	.w7(32'hbc5f1cf7),
	.w8(32'hbbb3d04b),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1e2ded),
	.w1(32'hbb9178c4),
	.w2(32'hbb10f73f),
	.w3(32'h3b8a63ba),
	.w4(32'hbbed8c9f),
	.w5(32'hbc03030f),
	.w6(32'hbb76db5d),
	.w7(32'h3b2930c6),
	.w8(32'hbb41d10e),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a95b9),
	.w1(32'hbb72ed54),
	.w2(32'hbb3cec42),
	.w3(32'hbbe40806),
	.w4(32'h3ce6f529),
	.w5(32'h3d27fb4d),
	.w6(32'hbb8e9972),
	.w7(32'hbcdb03a7),
	.w8(32'h3b1d5818),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba92816b),
	.w1(32'h3acb13a9),
	.w2(32'h3bf0abcd),
	.w3(32'h3caa5e65),
	.w4(32'h3c0bd061),
	.w5(32'h3c23b18a),
	.w6(32'hba35947a),
	.w7(32'hbc48daa8),
	.w8(32'hbb23bb48),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a982f95),
	.w1(32'hbb1ada8f),
	.w2(32'h3b49efa5),
	.w3(32'hb9945011),
	.w4(32'h3bb901ac),
	.w5(32'h3c3e0a05),
	.w6(32'hbc37b756),
	.w7(32'hbc6e3fa1),
	.w8(32'hbbb61c97),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0336ee),
	.w1(32'h3ab44799),
	.w2(32'h3c457a86),
	.w3(32'h3b8951d8),
	.w4(32'h3b4e5270),
	.w5(32'h3a5b2832),
	.w6(32'h3af99b2d),
	.w7(32'hbb9414f1),
	.w8(32'h3b077ae7),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb80893c),
	.w1(32'h3a8e2281),
	.w2(32'hbb850c77),
	.w3(32'hba219712),
	.w4(32'hb963ea5e),
	.w5(32'hbb127fa6),
	.w6(32'hbbe5b440),
	.w7(32'hbbff346c),
	.w8(32'hba9bcd07),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab38da2),
	.w1(32'hbba66fe3),
	.w2(32'hbb4a6de6),
	.w3(32'h3ad0b748),
	.w4(32'hbbf2e536),
	.w5(32'hbbeca211),
	.w6(32'hbb945fea),
	.w7(32'hb9d82f94),
	.w8(32'hbb9448fe),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba922e1),
	.w1(32'h3b9b3c5c),
	.w2(32'h3c242c02),
	.w3(32'hbbc91b8d),
	.w4(32'hbb31ad51),
	.w5(32'hbc0cdb62),
	.w6(32'h3c0e60d8),
	.w7(32'h3cac8b68),
	.w8(32'h3b441975),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1b670a),
	.w1(32'h3b373314),
	.w2(32'h3c1190cb),
	.w3(32'hbbc060c0),
	.w4(32'h3c031b3c),
	.w5(32'h3c548da6),
	.w6(32'hbb8dafab),
	.w7(32'hbc3fea27),
	.w8(32'hbb346130),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b03e1a2),
	.w1(32'hbbb740b4),
	.w2(32'h3c13bd1b),
	.w3(32'h3b472e0a),
	.w4(32'h3bceeebc),
	.w5(32'h3c5dca9f),
	.w6(32'hbb9ad68c),
	.w7(32'hbabd89a3),
	.w8(32'h3bf4bd84),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9dfb23),
	.w1(32'h3b96042f),
	.w2(32'h3b1df45a),
	.w3(32'hbbecc3f7),
	.w4(32'h3c138dfa),
	.w5(32'h3c443b6b),
	.w6(32'hbb316a40),
	.w7(32'hbb2855fb),
	.w8(32'hba987346),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb6bd89),
	.w1(32'hba0c186c),
	.w2(32'hbc014e05),
	.w3(32'h3c2fa4da),
	.w4(32'hb8d0854b),
	.w5(32'h3abe0085),
	.w6(32'h3b538dc2),
	.w7(32'hbc0800b2),
	.w8(32'hbbdd6200),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb097413),
	.w1(32'hbb6d3c38),
	.w2(32'hba158fb9),
	.w3(32'h3c6ef616),
	.w4(32'hb90e95e2),
	.w5(32'h3c0819cf),
	.w6(32'hbbef5b10),
	.w7(32'hbbdca0a1),
	.w8(32'hba899f84),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e9c280),
	.w1(32'hbbec6149),
	.w2(32'hbbf49589),
	.w3(32'h3b6eae0b),
	.w4(32'hbb1e9345),
	.w5(32'hba9e553c),
	.w6(32'hbbf37b75),
	.w7(32'hbaa79596),
	.w8(32'hb9c59867),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba905342),
	.w1(32'hbb6d96ed),
	.w2(32'h3b0fa52b),
	.w3(32'h3be080f0),
	.w4(32'h3a6c3ec4),
	.w5(32'h3c05ffb8),
	.w6(32'hbc010bbf),
	.w7(32'hbc24a82d),
	.w8(32'hbb0b055e),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be03eb4),
	.w1(32'h3aeb9421),
	.w2(32'h3b0961b5),
	.w3(32'h3bf937c9),
	.w4(32'hbb916cae),
	.w5(32'hbb7e36b6),
	.w6(32'h3a564698),
	.w7(32'h3b80829a),
	.w8(32'h3b922078),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb09fedc),
	.w1(32'hbbd8f89b),
	.w2(32'h3bb34b58),
	.w3(32'h3977f615),
	.w4(32'h3b7f88cb),
	.w5(32'h3c8a39c6),
	.w6(32'hbc8d2bc1),
	.w7(32'hbcb64719),
	.w8(32'hbc0b3695),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9fd8e4),
	.w1(32'hbbbb98d0),
	.w2(32'h3afddbb0),
	.w3(32'hb9628295),
	.w4(32'hbc1051eb),
	.w5(32'hbc1b6c92),
	.w6(32'hbab22a52),
	.w7(32'h3c515bca),
	.w8(32'hbaabb628),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb59eb7e),
	.w1(32'hbb834f6f),
	.w2(32'h3b35152f),
	.w3(32'hbba95ac6),
	.w4(32'h3955f786),
	.w5(32'h3c5ae62a),
	.w6(32'hbc4cb6b1),
	.w7(32'hbc906f32),
	.w8(32'hbc28a22c),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b49a6e9),
	.w1(32'hb96cf99d),
	.w2(32'h3bbf25db),
	.w3(32'h3b3aaa8a),
	.w4(32'hbbb593b8),
	.w5(32'hbc004f2a),
	.w6(32'h3a48377c),
	.w7(32'h3c3bdc22),
	.w8(32'h3b6e8eb5),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a65d0a0),
	.w1(32'hb9827c22),
	.w2(32'h3a98f4c5),
	.w3(32'hbb6c5482),
	.w4(32'h3c183f63),
	.w5(32'h3b904c3b),
	.w6(32'hbb4e3c34),
	.w7(32'hbb8b84fc),
	.w8(32'hbb612d1a),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c50bb13),
	.w1(32'hbb63e550),
	.w2(32'hbb46e0c2),
	.w3(32'h3c52f1ae),
	.w4(32'h3ca08167),
	.w5(32'h3cf916af),
	.w6(32'hbbc6605d),
	.w7(32'hbcb59535),
	.w8(32'hba113da3),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c6499a),
	.w1(32'hbb70c992),
	.w2(32'h3ad58e3f),
	.w3(32'h3c802ae3),
	.w4(32'h39301a56),
	.w5(32'h3c0e9698),
	.w6(32'hbc2ad912),
	.w7(32'hbc47d5d5),
	.w8(32'hbc2063bb),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acf487f),
	.w1(32'hbb2969d9),
	.w2(32'h3b79f503),
	.w3(32'h3b0344f0),
	.w4(32'hbbcb55f1),
	.w5(32'hbc059ece),
	.w6(32'h3aa8eb53),
	.w7(32'h3c089167),
	.w8(32'h3b99777c),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba361b8),
	.w1(32'hbb9cfb69),
	.w2(32'hbc0417af),
	.w3(32'hbbf96820),
	.w4(32'h3aa78d25),
	.w5(32'hba0c9998),
	.w6(32'hbbb80c5f),
	.w7(32'hbbd6b586),
	.w8(32'hba4f70b1),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b4cdb),
	.w1(32'hbbfaa870),
	.w2(32'hbc3ab2ef),
	.w3(32'h3bbcf0ea),
	.w4(32'hbb96395d),
	.w5(32'hbbd79fba),
	.w6(32'hbbd8977c),
	.w7(32'hbbf5ff03),
	.w8(32'hbb225316),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f597d),
	.w1(32'hbae6f7dc),
	.w2(32'h3b4e48fc),
	.w3(32'h3a641c0a),
	.w4(32'h3a1aa9a4),
	.w5(32'h39d1a16c),
	.w6(32'hbbba6f07),
	.w7(32'h3a85b666),
	.w8(32'hbb855588),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3193a0),
	.w1(32'h3bd39e58),
	.w2(32'h3c555143),
	.w3(32'h3aef8f14),
	.w4(32'h3b7e2c54),
	.w5(32'h3bae4a82),
	.w6(32'h3babf55d),
	.w7(32'h3be59820),
	.w8(32'h3a2e788b),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaffefb4),
	.w1(32'hbbaa5bbb),
	.w2(32'h3a052f35),
	.w3(32'hbb530575),
	.w4(32'h3c2ddc96),
	.w5(32'h3cc06b05),
	.w6(32'hbc708d9c),
	.w7(32'hbcd1df04),
	.w8(32'hbc1c4ac6),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa4ba67),
	.w1(32'hbbd54ae9),
	.w2(32'hba8d5fa9),
	.w3(32'h3c31d41a),
	.w4(32'hbbf17468),
	.w5(32'hbbf0bb90),
	.w6(32'hbb7f95b8),
	.w7(32'h3bd9c49f),
	.w8(32'hbbbf30bf),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe861b8),
	.w1(32'hbbb33c83),
	.w2(32'h3aa6d911),
	.w3(32'hbb606415),
	.w4(32'hbbc12113),
	.w5(32'hbbc248f1),
	.w6(32'hbb01f47d),
	.w7(32'h3c244e11),
	.w8(32'hba882959),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb17a99c),
	.w1(32'hbc33cd7f),
	.w2(32'hbc14841d),
	.w3(32'hbb28db24),
	.w4(32'hbbed27b0),
	.w5(32'hbbcf790f),
	.w6(32'hbc08941f),
	.w7(32'hbb0b22bc),
	.w8(32'hbc0744cf),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc19e904),
	.w1(32'hbb4ec322),
	.w2(32'h3b86f91d),
	.w3(32'hbb4eb08a),
	.w4(32'h3b6e18ea),
	.w5(32'h3c42ba36),
	.w6(32'hbc89aa80),
	.w7(32'hbca8ff1f),
	.w8(32'hbbe0e4c2),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b838618),
	.w1(32'h3a914c5f),
	.w2(32'h3c468543),
	.w3(32'hbb4cc866),
	.w4(32'hbbd121ef),
	.w5(32'h3ab7af10),
	.w6(32'h3c37737f),
	.w7(32'h3b402a0f),
	.w8(32'h3af07a37),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6e611b),
	.w1(32'hbb873e95),
	.w2(32'h39ef6faf),
	.w3(32'hbaaa37ef),
	.w4(32'hbc3c2a40),
	.w5(32'hbca53771),
	.w6(32'h3c235710),
	.w7(32'h3ce76309),
	.w8(32'h3b9811be),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc080c79),
	.w1(32'h3b15399b),
	.w2(32'h3c572329),
	.w3(32'hbc267b28),
	.w4(32'h3c07e53d),
	.w5(32'h3cb3c56f),
	.w6(32'hbbc8b4c7),
	.w7(32'hbc5648f1),
	.w8(32'hbb7f609d),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5100b4),
	.w1(32'h3b9d8011),
	.w2(32'h3c5f930c),
	.w3(32'h3c2164f7),
	.w4(32'hbac25852),
	.w5(32'hb995bb36),
	.w6(32'h3a8e1f1c),
	.w7(32'h3c137ba6),
	.w8(32'h3bbef49a),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab36ed3),
	.w1(32'hbc34ebb2),
	.w2(32'hbbc75449),
	.w3(32'hbb370427),
	.w4(32'hbc3a8bcf),
	.w5(32'hbc1fa7db),
	.w6(32'hbbd2f5e8),
	.w7(32'h3bc3695f),
	.w8(32'hbb607caf),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbfa75e),
	.w1(32'hbb92becb),
	.w2(32'hbc207e27),
	.w3(32'hbb832fde),
	.w4(32'hbb3ec030),
	.w5(32'hbb903b57),
	.w6(32'hbc084c71),
	.w7(32'hbc244f5e),
	.w8(32'hbb935e21),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1e59a1),
	.w1(32'hbb80dd2a),
	.w2(32'h3b197309),
	.w3(32'h3ace36fb),
	.w4(32'h384d9e94),
	.w5(32'h3c723781),
	.w6(32'hbc54d36b),
	.w7(32'hbca60fb9),
	.w8(32'hbc2541ba),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bece590),
	.w1(32'h3b677387),
	.w2(32'h3b44bb7f),
	.w3(32'h3c266935),
	.w4(32'h3b9db5c8),
	.w5(32'h3bbbf7d2),
	.w6(32'hbbd999c5),
	.w7(32'hbc047b13),
	.w8(32'hbae73f08),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39062b0d),
	.w1(32'hbbc1f2ad),
	.w2(32'h3aae120a),
	.w3(32'h3a0a73b4),
	.w4(32'h3b9dd685),
	.w5(32'h3c8634b0),
	.w6(32'hbc4d3ffe),
	.w7(32'hbc6c1df3),
	.w8(32'hbbbd9b43),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b483d29),
	.w1(32'h3b3fab6b),
	.w2(32'hbb7b59cd),
	.w3(32'h3b7d9ba6),
	.w4(32'hbbdac097),
	.w5(32'hbb20afc6),
	.w6(32'h3b293c11),
	.w7(32'hb8a3b490),
	.w8(32'hbbb780d8),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb19e240),
	.w1(32'hbac6766b),
	.w2(32'h3b4a990b),
	.w3(32'h39a54d6c),
	.w4(32'h3b24f242),
	.w5(32'h3bd9412d),
	.w6(32'hbbb6fce3),
	.w7(32'hbbe4dfa0),
	.w8(32'h3b387cb1),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b896123),
	.w1(32'hbb7c7f28),
	.w2(32'hba2620cc),
	.w3(32'h3b9ef315),
	.w4(32'hba42aa33),
	.w5(32'h39c86ba6),
	.w6(32'h3ac04a40),
	.w7(32'hbad572cd),
	.w8(32'hba8f44dc),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb810b76),
	.w1(32'hbc023ea4),
	.w2(32'hbbc1728b),
	.w3(32'hbb9cf886),
	.w4(32'hbbb60914),
	.w5(32'hbbadfb29),
	.w6(32'hbbbca220),
	.w7(32'h3aa5d24a),
	.w8(32'hbb58b1b5),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9e9b0b),
	.w1(32'h3a48fafc),
	.w2(32'h3aabfafe),
	.w3(32'hbb2adf6c),
	.w4(32'h3b90ecd0),
	.w5(32'h3c3b8ea9),
	.w6(32'hbb7e05c6),
	.w7(32'hbbf7acef),
	.w8(32'h3aae825b),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4d90d4),
	.w1(32'hbc2acf97),
	.w2(32'hbbe8ee9c),
	.w3(32'h3be3ba2d),
	.w4(32'hbc2dae0d),
	.w5(32'hbc2d40ac),
	.w6(32'hbbb9c427),
	.w7(32'h3baebd89),
	.w8(32'hbb1ef52b),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd2d627),
	.w1(32'hbc1e5483),
	.w2(32'hbc16360e),
	.w3(32'hbbb1f9d9),
	.w4(32'hbbcb35a3),
	.w5(32'hbbe27073),
	.w6(32'hbbedc7cb),
	.w7(32'hbabb89a0),
	.w8(32'hbbf21e9f),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc098d37),
	.w1(32'hbae50dc0),
	.w2(32'hbb47a143),
	.w3(32'hbb8bf0b8),
	.w4(32'h3c0ef288),
	.w5(32'h3c97048b),
	.w6(32'hbc117773),
	.w7(32'hbcba6ac8),
	.w8(32'hbbd81f52),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3bb7d0),
	.w1(32'hbb3c3baf),
	.w2(32'hbb8926a5),
	.w3(32'h3c340c29),
	.w4(32'h3c3f2dfb),
	.w5(32'h3cb11dac),
	.w6(32'hbc428640),
	.w7(32'hbc8c621f),
	.w8(32'hbbd103c7),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b833be9),
	.w1(32'hbc13165e),
	.w2(32'hbc352171),
	.w3(32'h3c688f56),
	.w4(32'hbbb2a6e2),
	.w5(32'hbb992536),
	.w6(32'hbc5323a2),
	.w7(32'hbc382e6f),
	.w8(32'hbba0b611),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac59bf4),
	.w1(32'hbc39483f),
	.w2(32'hbc32a3ca),
	.w3(32'h3b10bec6),
	.w4(32'hbb0eee25),
	.w5(32'h3b6bd432),
	.w6(32'hbc141ec7),
	.w7(32'hbc5920b3),
	.w8(32'hbbc08043),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc02a430),
	.w1(32'hbc021320),
	.w2(32'hbbde9dfa),
	.w3(32'h38f30543),
	.w4(32'hb8cc4edf),
	.w5(32'h39e67448),
	.w6(32'hbbaec54b),
	.w7(32'hbc05425a),
	.w8(32'hbc6d793a),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0cec0a),
	.w1(32'h3b485719),
	.w2(32'h3b2d9a9e),
	.w3(32'h3c403606),
	.w4(32'hb98c603f),
	.w5(32'h3abd473f),
	.w6(32'h3b3a8866),
	.w7(32'hba1969ce),
	.w8(32'hbb88923c),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba810b0d),
	.w1(32'hbbe3b550),
	.w2(32'hbb243009),
	.w3(32'hba52b9b2),
	.w4(32'h3ad70a56),
	.w5(32'h3b94c800),
	.w6(32'hbbbe62d4),
	.w7(32'h3bb19a1e),
	.w8(32'h3adfeb8d),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e211e),
	.w1(32'hbbcefd3b),
	.w2(32'hba48b50f),
	.w3(32'hbc0b6b94),
	.w4(32'hbabc8d5f),
	.w5(32'h3c8a2bba),
	.w6(32'hbca1ee20),
	.w7(32'hbceb2e82),
	.w8(32'hbc8b5be3),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb4b0e5),
	.w1(32'hbb36ad12),
	.w2(32'hba6cecbb),
	.w3(32'h3c55d6a4),
	.w4(32'h3bb1c59d),
	.w5(32'h3c756d9c),
	.w6(32'hbc0c4c76),
	.w7(32'hbc525a67),
	.w8(32'h3a48c978),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb49308),
	.w1(32'h3b6e9c45),
	.w2(32'h3c4dc559),
	.w3(32'h3c33e760),
	.w4(32'hbb19b183),
	.w5(32'h3b83dce7),
	.w6(32'hbb04169a),
	.w7(32'hbb82b31a),
	.w8(32'hbac132c3),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd7bfa8),
	.w1(32'h3a758ede),
	.w2(32'h3beacca4),
	.w3(32'h3bbe9d22),
	.w4(32'hbc1d7b3e),
	.w5(32'hbc8982ea),
	.w6(32'h3bbea63b),
	.w7(32'hba5b6a7d),
	.w8(32'hbb7315d6),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbda3aa2),
	.w1(32'hbbca87a0),
	.w2(32'h3a5cb9fb),
	.w3(32'h3c173aa3),
	.w4(32'hbc900615),
	.w5(32'hbcff837d),
	.w6(32'h3c793229),
	.w7(32'h3d2f9033),
	.w8(32'h3beed692),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4e4aa7),
	.w1(32'hbbce1e2a),
	.w2(32'hba46df65),
	.w3(32'hbc81de7b),
	.w4(32'hbbeea467),
	.w5(32'hbbc8c30f),
	.w6(32'hbb8cad99),
	.w7(32'h3bdd3656),
	.w8(32'hbbe99451),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcba587),
	.w1(32'hbb4e873c),
	.w2(32'hb65deb3e),
	.w3(32'hbaef65b9),
	.w4(32'hbc0175a1),
	.w5(32'hbc64c1d0),
	.w6(32'h3bede64c),
	.w7(32'h3cac0dc4),
	.w8(32'h3b5ec0be),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc5bc87),
	.w1(32'hbb377908),
	.w2(32'hb9b2c11a),
	.w3(32'hbbda6337),
	.w4(32'hbbbcad3d),
	.w5(32'hbbb07b87),
	.w6(32'hbaf9e481),
	.w7(32'h3b930da2),
	.w8(32'h3a3c243f),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e23ad8),
	.w1(32'hbc76ba9d),
	.w2(32'hbc09ec0a),
	.w3(32'hbb18bcf9),
	.w4(32'h39b57bf3),
	.w5(32'h3be6c94f),
	.w6(32'hbc4646d2),
	.w7(32'hbc5927ba),
	.w8(32'hbb0da25d),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad58eb7),
	.w1(32'hbc5a56cc),
	.w2(32'hbc401580),
	.w3(32'h3bc14605),
	.w4(32'hbbce5a74),
	.w5(32'hbbe959cd),
	.w6(32'hbc11546f),
	.w7(32'hb9301289),
	.w8(32'hbbd9e1e0),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc29b557),
	.w1(32'hbb5a6905),
	.w2(32'h39ff8116),
	.w3(32'hbb7d97bf),
	.w4(32'hbc1f304e),
	.w5(32'hbc8caa09),
	.w6(32'h3bff028f),
	.w7(32'h3cb753b0),
	.w8(32'h3b5db80a),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdf8b43),
	.w1(32'hb9045e72),
	.w2(32'h3bd1d005),
	.w3(32'hbc11e725),
	.w4(32'h3c076224),
	.w5(32'h3c90e683),
	.w6(32'hbbb8cf92),
	.w7(32'hbc949a51),
	.w8(32'hbc4dee46),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a20b352),
	.w1(32'hbb9e2ece),
	.w2(32'h3abfb270),
	.w3(32'h3c15c574),
	.w4(32'hba0b41ac),
	.w5(32'h3b0ce783),
	.w6(32'hbc080b30),
	.w7(32'h3b26f17f),
	.w8(32'hbab9c2be),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b289d89),
	.w1(32'hba7f6d8f),
	.w2(32'hbaae804f),
	.w3(32'h3b18e501),
	.w4(32'h3ae72c77),
	.w5(32'h3b60dd86),
	.w6(32'h3c16e7ee),
	.w7(32'h3b8da480),
	.w8(32'hbab2ea21),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a56eb9d),
	.w1(32'hbb37da75),
	.w2(32'h3b3879ab),
	.w3(32'hbab867db),
	.w4(32'h3b03ad2c),
	.w5(32'h3b7f84ef),
	.w6(32'hbbbdde3f),
	.w7(32'h3a949d18),
	.w8(32'h3a138f0d),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1dbd30),
	.w1(32'hbb750d1e),
	.w2(32'h3b94c908),
	.w3(32'h3b6386ff),
	.w4(32'h3b8e3f15),
	.w5(32'h3c4e8ad8),
	.w6(32'hbbfbdc3f),
	.w7(32'hbc25bf3b),
	.w8(32'hb94cec21),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b448086),
	.w1(32'hbabc8362),
	.w2(32'h3b3fbcb3),
	.w3(32'h3b85b702),
	.w4(32'hbbd34fcf),
	.w5(32'hbbf776eb),
	.w6(32'hbb92b4a2),
	.w7(32'h3b8c2b83),
	.w8(32'hbbaa2616),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb93d652),
	.w1(32'hbb976c17),
	.w2(32'h3a02299d),
	.w3(32'hbbcf0272),
	.w4(32'hbc541b05),
	.w5(32'hbcbb3ce8),
	.w6(32'h3c394cfb),
	.w7(32'h3d03248f),
	.w8(32'h3baa26be),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1a4d6c),
	.w1(32'hb98599cf),
	.w2(32'h3b7a8326),
	.w3(32'hbc3c7912),
	.w4(32'hbba07136),
	.w5(32'hbbf9ddcf),
	.w6(32'h3b95b7f8),
	.w7(32'h3c8b0dc1),
	.w8(32'h3b359988),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaca1edd),
	.w1(32'hb994e568),
	.w2(32'h3acd9ee7),
	.w3(32'hbafd7e2c),
	.w4(32'hbb8ccafb),
	.w5(32'hbbe49247),
	.w6(32'h3ba7b117),
	.w7(32'h3c883ec0),
	.w8(32'h3b45d6b5),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba61e1f2),
	.w1(32'hbbc9d433),
	.w2(32'hba2452a0),
	.w3(32'h3a22b118),
	.w4(32'hbc253645),
	.w5(32'hbc9e0ac8),
	.w6(32'hbbc0ab7e),
	.w7(32'h39a5b705),
	.w8(32'hba5c03c0),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc220c17),
	.w1(32'h3b843a15),
	.w2(32'h3c1fba7a),
	.w3(32'hbc20e59b),
	.w4(32'h3b947d86),
	.w5(32'h3c712429),
	.w6(32'hbbab45c6),
	.w7(32'hbc0ea3be),
	.w8(32'hb8ebbdee),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39fc9c45),
	.w1(32'hbb33e063),
	.w2(32'hbb8720b8),
	.w3(32'h3b2bb390),
	.w4(32'hb9fa9541),
	.w5(32'h3b358fdc),
	.w6(32'hbbb9a68c),
	.w7(32'hbb9036fe),
	.w8(32'hbc13f5ec),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba40c5d5),
	.w1(32'hba661059),
	.w2(32'hba2365fc),
	.w3(32'h3bcddfaf),
	.w4(32'h3b596dea),
	.w5(32'h3baa5d16),
	.w6(32'hbb72f86d),
	.w7(32'hbb8ccbad),
	.w8(32'hbaf2e7fa),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a251f1a),
	.w1(32'hbb2eb18c),
	.w2(32'h3b9b261f),
	.w3(32'h3b9bd1e6),
	.w4(32'hbc058ddd),
	.w5(32'hbc2268c4),
	.w6(32'h3b173ac0),
	.w7(32'h3c8b83ef),
	.w8(32'hb941d0e8),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4f974b),
	.w1(32'hbb506325),
	.w2(32'h3c3ad64c),
	.w3(32'hbbbeb673),
	.w4(32'hbbaf2449),
	.w5(32'hbc349c53),
	.w6(32'hbb773e23),
	.w7(32'hbb404cca),
	.w8(32'hbbbb571a),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb48858e),
	.w1(32'hb9aed1ce),
	.w2(32'hba8e2d0f),
	.w3(32'h3923015b),
	.w4(32'h3bb2fe9f),
	.w5(32'h3c3aa69d),
	.w6(32'hbbdd85b3),
	.w7(32'hbc2e4027),
	.w8(32'hbc482c7a),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b11b0cd),
	.w1(32'hbc517902),
	.w2(32'hbc09a93c),
	.w3(32'h3c79f87d),
	.w4(32'hbc1a982f),
	.w5(32'hbbf8bc02),
	.w6(32'hbc1960b9),
	.w7(32'hba12004b),
	.w8(32'hbbcb2c1f),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd30c64),
	.w1(32'hb66347a6),
	.w2(32'h3682941e),
	.w3(32'hbb512a3d),
	.w4(32'hb60ce416),
	.w5(32'h36a51322),
	.w6(32'h360d4514),
	.w7(32'h367caf85),
	.w8(32'h372a3d35),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6f45e98),
	.w1(32'hb800aea4),
	.w2(32'hb7af044d),
	.w3(32'h37f26f74),
	.w4(32'h34dbfa0f),
	.w5(32'h36c706a9),
	.w6(32'h380456f5),
	.w7(32'h37d0a44c),
	.w8(32'h36a30d05),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule