module layer_10_featuremap_335(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb306b2b),
	.w1(32'hb81a79be),
	.w2(32'h3b2b056b),
	.w3(32'h3b301916),
	.w4(32'h3bc378c9),
	.w5(32'hbb98c57e),
	.w6(32'h3a6e2e3d),
	.w7(32'h3b944d80),
	.w8(32'hbb6f60be),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7964e9),
	.w1(32'hbb3aa1c0),
	.w2(32'hbaf2ce1e),
	.w3(32'hbbba4893),
	.w4(32'hbb80b4b3),
	.w5(32'h3bd29bf7),
	.w6(32'hbb87801c),
	.w7(32'hba9d140e),
	.w8(32'h3c01b08d),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b02e2cb),
	.w1(32'hba838c3c),
	.w2(32'hbadfceaa),
	.w3(32'h3bbeef43),
	.w4(32'h3b899691),
	.w5(32'h3b12546d),
	.w6(32'h3ba0e9e6),
	.w7(32'h3b3a0f22),
	.w8(32'h3b2a679a),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2ce456),
	.w1(32'h3b0224e6),
	.w2(32'h3a8dee59),
	.w3(32'h3a1168d0),
	.w4(32'hba89d644),
	.w5(32'h3b7fc125),
	.w6(32'h3a614e70),
	.w7(32'hba197699),
	.w8(32'hbb45614b),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be8e827),
	.w1(32'h3c0010bc),
	.w2(32'h3c53644b),
	.w3(32'h3bb0551a),
	.w4(32'h3c26700a),
	.w5(32'h3b72782c),
	.w6(32'hbb729d25),
	.w7(32'h3b7ab168),
	.w8(32'h3ad8e45f),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1d39c9),
	.w1(32'h3af07de8),
	.w2(32'h3a1e3e3b),
	.w3(32'h3b0873bc),
	.w4(32'h3a9d095d),
	.w5(32'h3b7fb54c),
	.w6(32'hb84f6c2c),
	.w7(32'hb997c85d),
	.w8(32'h3bb24b67),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bce461f),
	.w1(32'h3b8c2ea4),
	.w2(32'h3b549cd8),
	.w3(32'h3afdae87),
	.w4(32'h391edc55),
	.w5(32'hb917c003),
	.w6(32'h3b674170),
	.w7(32'h3aa20ed4),
	.w8(32'h3a34c73f),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b2dce5),
	.w1(32'h3a5ce2e9),
	.w2(32'h39122b23),
	.w3(32'h3b82e280),
	.w4(32'h3afa5742),
	.w5(32'h3bb53eb3),
	.w6(32'h3b52b3e9),
	.w7(32'h39a04a5c),
	.w8(32'h3b9c34f0),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7c51cf),
	.w1(32'h3b598b5a),
	.w2(32'h3a88ff9f),
	.w3(32'h3b7e62e2),
	.w4(32'h3b1146b5),
	.w5(32'h3b8188c5),
	.w6(32'h3b52c320),
	.w7(32'h39d4916c),
	.w8(32'h3a84abff),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a589f79),
	.w1(32'h39bfdf29),
	.w2(32'h3a02a6b8),
	.w3(32'hb88701b8),
	.w4(32'hba75ea14),
	.w5(32'h3b9ccd44),
	.w6(32'hbb29b0bf),
	.w7(32'hbb44ae23),
	.w8(32'h3afdee4b),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaaa2e9),
	.w1(32'h3b06f143),
	.w2(32'h3b5df8d2),
	.w3(32'h3ac390fd),
	.w4(32'h3b452dd4),
	.w5(32'hbb666799),
	.w6(32'hba9d8d45),
	.w7(32'h3ac5ba71),
	.w8(32'hb9457b76),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a30db2a),
	.w1(32'hba176088),
	.w2(32'hba29a8d5),
	.w3(32'hba65fd95),
	.w4(32'hba7c2879),
	.w5(32'hbb4b3b75),
	.w6(32'h3afbae9e),
	.w7(32'h3ab688d9),
	.w8(32'hbafd1db4),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb01e896),
	.w1(32'hb969f654),
	.w2(32'h3bbcebe9),
	.w3(32'hbb903a6e),
	.w4(32'h38d19efa),
	.w5(32'hbab1c154),
	.w6(32'hbb8bf19e),
	.w7(32'hbae2e05c),
	.w8(32'hbb1f7f4f),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb172a84),
	.w1(32'h3ac0fc3d),
	.w2(32'h3bc0f245),
	.w3(32'hb5ee9bf5),
	.w4(32'h3bad8d52),
	.w5(32'h3b84c692),
	.w6(32'hbab5c648),
	.w7(32'h3b9a8cce),
	.w8(32'h3b8b530d),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b549130),
	.w1(32'h3b22c33a),
	.w2(32'h3b351a4e),
	.w3(32'h3b574356),
	.w4(32'h3b1a750d),
	.w5(32'hb93c31f7),
	.w6(32'h3b600c61),
	.w7(32'hb95eba46),
	.w8(32'hbb00a5b3),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa5442c),
	.w1(32'hbb742a52),
	.w2(32'hbb3ddf5f),
	.w3(32'hbba31435),
	.w4(32'hbb689d93),
	.w5(32'h3be2e836),
	.w6(32'hbba923e0),
	.w7(32'hbb222b29),
	.w8(32'h3bd31e44),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b841358),
	.w1(32'h3b4362b4),
	.w2(32'h3b210ebd),
	.w3(32'h3b9fd48c),
	.w4(32'h3ad28170),
	.w5(32'hb8ab39f5),
	.w6(32'h3b81fed5),
	.w7(32'h3a5876dd),
	.w8(32'hba449e6e),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba618e3d),
	.w1(32'hba2283d8),
	.w2(32'h3b5d3741),
	.w3(32'h3ad0c454),
	.w4(32'h3a91420d),
	.w5(32'h3afb3229),
	.w6(32'h3aee9115),
	.w7(32'h3ad89047),
	.w8(32'h3b227c7e),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafa45a4),
	.w1(32'hbaa83dae),
	.w2(32'h3ab1e5fa),
	.w3(32'h3986d1f5),
	.w4(32'h3ab694f0),
	.w5(32'h38b5185f),
	.w6(32'hbae055db),
	.w7(32'hbb0f87e9),
	.w8(32'h3bbfb3fa),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c032d79),
	.w1(32'h3b934b4d),
	.w2(32'h3b048c88),
	.w3(32'hbbc3563c),
	.w4(32'hbb916b36),
	.w5(32'h3b20b20b),
	.w6(32'hbb500028),
	.w7(32'hbb859ba7),
	.w8(32'h3b1c44ea),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b87b0f6),
	.w1(32'hbb0f8220),
	.w2(32'hbb6f7389),
	.w3(32'hbb40239e),
	.w4(32'hbb7b8d3d),
	.w5(32'h3b57dd5c),
	.w6(32'hbb3f8f08),
	.w7(32'hbb5537db),
	.w8(32'h3b844cb2),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6be83a),
	.w1(32'h3b80a33b),
	.w2(32'h3b4ea419),
	.w3(32'h3b29589f),
	.w4(32'h3ac58b3e),
	.w5(32'hbb647539),
	.w6(32'h3b96860d),
	.w7(32'h3b30c232),
	.w8(32'hbbb156c9),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e36fd6),
	.w1(32'h3a9e41f9),
	.w2(32'hba6edfb4),
	.w3(32'hbb0afb8b),
	.w4(32'h38cf6a8d),
	.w5(32'hb89f8197),
	.w6(32'hb9b491e4),
	.w7(32'h3b5c142d),
	.w8(32'h39317732),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7bf828),
	.w1(32'hbb9411d1),
	.w2(32'hbb1b157c),
	.w3(32'hbbf23aec),
	.w4(32'hbb4da3d3),
	.w5(32'h3b97915d),
	.w6(32'hbc091cae),
	.w7(32'hbae1fbd5),
	.w8(32'h3a672937),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf9cef6),
	.w1(32'hbbf0b181),
	.w2(32'hbb904e26),
	.w3(32'h3b2653cd),
	.w4(32'hb99308f2),
	.w5(32'h3b4004bf),
	.w6(32'hbaf6a3d1),
	.w7(32'hba203369),
	.w8(32'h3ba5f7e7),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b610767),
	.w1(32'h3b541773),
	.w2(32'hb7a36d9a),
	.w3(32'h3ad8f843),
	.w4(32'h3a093be2),
	.w5(32'h3b470e49),
	.w6(32'h3b87034a),
	.w7(32'hb79535c9),
	.w8(32'h3b1f12a5),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acbeb75),
	.w1(32'h3b66e1a2),
	.w2(32'h3b99128e),
	.w3(32'h3bc9d392),
	.w4(32'h3c03612e),
	.w5(32'hb60030d3),
	.w6(32'h3bacba7c),
	.w7(32'h3bcd568e),
	.w8(32'hbb5fb49d),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb83264f),
	.w1(32'hbba50dac),
	.w2(32'hbb909135),
	.w3(32'hbb071988),
	.w4(32'hbae5ee2d),
	.w5(32'h3a497d98),
	.w6(32'hbbae2064),
	.w7(32'hbba1c6cc),
	.w8(32'hbb97d250),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc27e5a),
	.w1(32'hbb3943f6),
	.w2(32'h3a6f313c),
	.w3(32'h3bfe23f5),
	.w4(32'h3c0f8c48),
	.w5(32'h3afb411b),
	.w6(32'h3aced236),
	.w7(32'h3bc0c752),
	.w8(32'h3b2f9506),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8961b8),
	.w1(32'h3ad41146),
	.w2(32'h3bafb26a),
	.w3(32'hbb171c0c),
	.w4(32'h3b593fef),
	.w5(32'h3b01b3f6),
	.w6(32'hbb7b75ef),
	.w7(32'h3b61178d),
	.w8(32'h3b9db2a8),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4efc58),
	.w1(32'h3c860ea6),
	.w2(32'h3c44a2ca),
	.w3(32'h3b31dbe6),
	.w4(32'h3bb93b89),
	.w5(32'h3c1964e9),
	.w6(32'h3b815f92),
	.w7(32'h3bd373cc),
	.w8(32'h3c124433),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb993a208),
	.w1(32'hba07027f),
	.w2(32'h3a8e9434),
	.w3(32'h3c13b4a9),
	.w4(32'h3bd4a0c1),
	.w5(32'hbb33e442),
	.w6(32'h3c0015a5),
	.w7(32'h3bec30eb),
	.w8(32'hbb597131),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb763ea1),
	.w1(32'hbbbcb8c8),
	.w2(32'hbc037849),
	.w3(32'hbaba3c01),
	.w4(32'hba923a48),
	.w5(32'h39eacc4b),
	.w6(32'hbb3e9b33),
	.w7(32'hbba6d64a),
	.w8(32'hb911aae0),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2f881b),
	.w1(32'hbb094889),
	.w2(32'h3a12c183),
	.w3(32'hba9b9f5a),
	.w4(32'h3a031aec),
	.w5(32'h3bfd4c75),
	.w6(32'hbb06c347),
	.w7(32'hb9c96c3b),
	.w8(32'h3b0f7b09),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9221284),
	.w1(32'hbaf1c575),
	.w2(32'h3b70aa63),
	.w3(32'h3c15bba8),
	.w4(32'h3bf678d7),
	.w5(32'h3b98dcf0),
	.w6(32'h3b9a03e2),
	.w7(32'h3c1b13a1),
	.w8(32'h3b7ee713),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad706a4),
	.w1(32'hba3fdb37),
	.w2(32'h3a8d3299),
	.w3(32'h3b7aefea),
	.w4(32'h3b2aa4d1),
	.w5(32'h3a1282a8),
	.w6(32'h3b6ecf76),
	.w7(32'h3a925535),
	.w8(32'hb93571ae),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a19c4a4),
	.w1(32'h3a7832ae),
	.w2(32'hba1f4395),
	.w3(32'h3a8b956c),
	.w4(32'h39abcfd0),
	.w5(32'hbaf9966b),
	.w6(32'h3b2d70d1),
	.w7(32'h3ab80300),
	.w8(32'hba6d8a0f),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a315747),
	.w1(32'hb9ff0109),
	.w2(32'hbb85964a),
	.w3(32'hbb0a2a26),
	.w4(32'hba4b1f9c),
	.w5(32'h3b0c6677),
	.w6(32'hbabfef17),
	.w7(32'hbb04072f),
	.w8(32'hbb3d1de6),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb856be9),
	.w1(32'hbba200f1),
	.w2(32'hbb9e3de0),
	.w3(32'h3a3bd6b1),
	.w4(32'h3aaf1ddb),
	.w5(32'h3aac3df6),
	.w6(32'hbb817172),
	.w7(32'hba625098),
	.w8(32'hb9838218),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1b2bce),
	.w1(32'h3aa2fdf6),
	.w2(32'h3b7c3d11),
	.w3(32'hbae88df1),
	.w4(32'hba802913),
	.w5(32'hbb72eb8a),
	.w6(32'hbad6423e),
	.w7(32'h3a77d58a),
	.w8(32'hbb9831c2),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6d8718),
	.w1(32'h3b1534f5),
	.w2(32'h3b8efd35),
	.w3(32'h3881d770),
	.w4(32'h3b639898),
	.w5(32'h3ab0d5c4),
	.w6(32'h3aaca53d),
	.w7(32'h3bd64cbb),
	.w8(32'h3aedcbf6),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d75697),
	.w1(32'hb9603883),
	.w2(32'hba8e0b3e),
	.w3(32'hb9833b4e),
	.w4(32'hba20ac5a),
	.w5(32'h38f2f68f),
	.w6(32'h3a866dbc),
	.w7(32'hba841ef0),
	.w8(32'hbaef6c62),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390c30ae),
	.w1(32'hbabf30d3),
	.w2(32'hba723707),
	.w3(32'h3941f055),
	.w4(32'h3a9b2751),
	.w5(32'hbb3aaae8),
	.w6(32'hbab8c0cc),
	.w7(32'hbad32781),
	.w8(32'hbb76a6e5),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9f714b),
	.w1(32'hb9f5b43d),
	.w2(32'h3b074e65),
	.w3(32'hbb83f850),
	.w4(32'hbb012c0f),
	.w5(32'h3bd11a33),
	.w6(32'hbb24b65e),
	.w7(32'hba91d1a1),
	.w8(32'h3c05bd8f),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b676325),
	.w1(32'h3bad4450),
	.w2(32'h3b75a8d8),
	.w3(32'h3b7506cf),
	.w4(32'h3b40db5d),
	.w5(32'hbb0f366e),
	.w6(32'h3bc92207),
	.w7(32'h3b81a5c8),
	.w8(32'hbb360c80),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba90d53d),
	.w1(32'h3aba9520),
	.w2(32'h3a4faf9f),
	.w3(32'hbb2294b3),
	.w4(32'hba3b4a72),
	.w5(32'h38c1fb2c),
	.w6(32'hbb725b5c),
	.w7(32'hbad0e748),
	.w8(32'hbaba5262),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2026d0),
	.w1(32'hbaa2c391),
	.w2(32'hbb043fb8),
	.w3(32'hbaae045e),
	.w4(32'hba7e1154),
	.w5(32'h3b9e148a),
	.w6(32'hbab7bff7),
	.w7(32'hbad58dd6),
	.w8(32'h3bb0489e),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8514ad),
	.w1(32'h3b24b373),
	.w2(32'h3b307b76),
	.w3(32'h3ba69293),
	.w4(32'hba81c656),
	.w5(32'h39a58e6e),
	.w6(32'h3bdad91c),
	.w7(32'h3a5572e2),
	.w8(32'h3a6065b0),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadce330),
	.w1(32'hbad322c7),
	.w2(32'hbade9e19),
	.w3(32'hba88e4b9),
	.w4(32'hb9acafdf),
	.w5(32'h3b584351),
	.w6(32'hba87ad10),
	.w7(32'hbae656e1),
	.w8(32'h3b6f75af),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6dc695),
	.w1(32'h3b88878b),
	.w2(32'h3b47fba8),
	.w3(32'h3b4435c1),
	.w4(32'h3ad048a0),
	.w5(32'hbb93174c),
	.w6(32'h3b8a696e),
	.w7(32'h3ad48f70),
	.w8(32'hbb4c6c23),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb745292),
	.w1(32'hb9c5bbb1),
	.w2(32'h3b69c1a9),
	.w3(32'hba964965),
	.w4(32'h3b4b01f1),
	.w5(32'hbacf4851),
	.w6(32'hba9b5f2e),
	.w7(32'h3b026f8f),
	.w8(32'hba20c1c5),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb182634),
	.w1(32'hb9a51c2c),
	.w2(32'h3a3eada6),
	.w3(32'hbb36ff5e),
	.w4(32'hbacc7f58),
	.w5(32'hbb65dd7a),
	.w6(32'hbb5d5645),
	.w7(32'hbab49edf),
	.w8(32'hbb3887b8),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbaef12),
	.w1(32'hbad14281),
	.w2(32'h39e739e4),
	.w3(32'hbb027120),
	.w4(32'h39d03398),
	.w5(32'h3b8ad2d5),
	.w6(32'hbac9f567),
	.w7(32'h3ad4fcbb),
	.w8(32'h3b1fef89),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b714686),
	.w1(32'h3c183457),
	.w2(32'h3c0dbeac),
	.w3(32'h3bc6a662),
	.w4(32'h3b9c3e7b),
	.w5(32'hbaccb078),
	.w6(32'h3bb6e832),
	.w7(32'h3bba9905),
	.w8(32'h3b98051e),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baf9658),
	.w1(32'h3b4e40ea),
	.w2(32'hb9a731c1),
	.w3(32'hbbdf6cc9),
	.w4(32'hbc14a4c3),
	.w5(32'h3b3722b2),
	.w6(32'hbb595ea0),
	.w7(32'hbbb8be0c),
	.w8(32'h39c30d96),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8a61e1),
	.w1(32'h395fcab7),
	.w2(32'h3bda413e),
	.w3(32'h3bc4e1ac),
	.w4(32'h3bb1230d),
	.w5(32'hba0a5629),
	.w6(32'h3b8efd63),
	.w7(32'h3c1ed053),
	.w8(32'hbab437cc),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb08527e),
	.w1(32'h3b164196),
	.w2(32'h3be9ec76),
	.w3(32'h3ba064d4),
	.w4(32'h3ba9ec23),
	.w5(32'h3c10f5ce),
	.w6(32'h3bd5da81),
	.w7(32'h3c37bc41),
	.w8(32'h3c28829f),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c14fda5),
	.w1(32'h3b599a99),
	.w2(32'hb9c4d15d),
	.w3(32'h3a96d208),
	.w4(32'hba8df55b),
	.w5(32'h3b642e4d),
	.w6(32'hbaadf423),
	.w7(32'hba9c9ba8),
	.w8(32'h3b9d0253),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b867a2d),
	.w1(32'h3b801ebb),
	.w2(32'h3b46ac62),
	.w3(32'h3b548686),
	.w4(32'h3af446a9),
	.w5(32'hb6118655),
	.w6(32'h3bb9fdfb),
	.w7(32'h3b1dd17a),
	.w8(32'h3b586b90),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b047704),
	.w1(32'h3b038f62),
	.w2(32'h39665c90),
	.w3(32'h3b247462),
	.w4(32'h39c7a27d),
	.w5(32'hba0943da),
	.w6(32'h3b85f4bc),
	.w7(32'h3aa440d2),
	.w8(32'hbb21cb2c),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb273095),
	.w1(32'hbb05ac4b),
	.w2(32'hbae7215a),
	.w3(32'hbaa6d5a1),
	.w4(32'hba85dc46),
	.w5(32'hbb0ede3b),
	.w6(32'hbb627d9b),
	.w7(32'hbb52803e),
	.w8(32'h3a43227a),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97de581),
	.w1(32'h397f96c9),
	.w2(32'hbad48ae7),
	.w3(32'hbb1acb77),
	.w4(32'hbb19add9),
	.w5(32'h3b090f9c),
	.w6(32'hba5e1de4),
	.w7(32'hbab6d057),
	.w8(32'hbacecd8d),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb50b1a9),
	.w1(32'hbb6c6821),
	.w2(32'hbaccffbc),
	.w3(32'h3b4e124a),
	.w4(32'h3b08e6dd),
	.w5(32'hbb020708),
	.w6(32'hbb067bfc),
	.w7(32'h3a0a2c57),
	.w8(32'hbb3de5bc),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2929e2),
	.w1(32'hba779fd3),
	.w2(32'h3b892b15),
	.w3(32'h39eda9b8),
	.w4(32'h3b4665ae),
	.w5(32'hbae0b2cb),
	.w6(32'h3a5cdc76),
	.w7(32'h3bed5bc7),
	.w8(32'hb9ae53ec),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb728626a),
	.w1(32'hbb02d7af),
	.w2(32'h3b34ea41),
	.w3(32'h39b20da0),
	.w4(32'h3ae182ef),
	.w5(32'hbbd4fdd7),
	.w6(32'hba78f30b),
	.w7(32'h3bf08d43),
	.w8(32'hbb4f4586),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5f3225),
	.w1(32'h3ba5f993),
	.w2(32'h3b55308a),
	.w3(32'hbbecc0e1),
	.w4(32'hbbd4567d),
	.w5(32'h3b8ad8b0),
	.w6(32'hbb88c51d),
	.w7(32'hbb732353),
	.w8(32'h3b49fb7b),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9d4243),
	.w1(32'hbb362a8d),
	.w2(32'hbafa9219),
	.w3(32'h3ae50da7),
	.w4(32'hba77a4a7),
	.w5(32'h3a64c9f3),
	.w6(32'hb9aba1ce),
	.w7(32'hbb577dcf),
	.w8(32'h3a798c14),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba395d20),
	.w1(32'h3a6d6a1e),
	.w2(32'h3b2abc43),
	.w3(32'h3aa26706),
	.w4(32'h3a67b388),
	.w5(32'hbaedef67),
	.w6(32'h3b08f140),
	.w7(32'h3a688753),
	.w8(32'h3993f5d5),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae445a0),
	.w1(32'hbbeeff6a),
	.w2(32'hbbe22f0d),
	.w3(32'hbbde57b6),
	.w4(32'hbbe799ba),
	.w5(32'h3b547596),
	.w6(32'hbbb9c845),
	.w7(32'hbb8471b1),
	.w8(32'h3b284e09),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ea0eda),
	.w1(32'h3a71cc43),
	.w2(32'h3bd5d4e9),
	.w3(32'hb89e9903),
	.w4(32'h3b1a4e5e),
	.w5(32'h3ae4deb8),
	.w6(32'hb9d04cb7),
	.w7(32'h399ee8d7),
	.w8(32'h3a400605),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d23594),
	.w1(32'h398d76dd),
	.w2(32'hbae72d3b),
	.w3(32'h3992f593),
	.w4(32'hb9e20d78),
	.w5(32'h3b03bac6),
	.w6(32'h3a1adad0),
	.w7(32'hbaf7c65d),
	.w8(32'h39b09bd5),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab47682),
	.w1(32'h396fbf58),
	.w2(32'h3a18b702),
	.w3(32'hb9177e2c),
	.w4(32'hbaac7110),
	.w5(32'hb9ca3b11),
	.w6(32'hbae5555a),
	.w7(32'hb9e42c9e),
	.w8(32'h3b00d7bd),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb527c81),
	.w1(32'hbb51b469),
	.w2(32'hbb604c9d),
	.w3(32'hbabe5950),
	.w4(32'hbb1f8414),
	.w5(32'hba079a96),
	.w6(32'h3a42a286),
	.w7(32'hb83c1f54),
	.w8(32'hba213d59),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4a7c34),
	.w1(32'hb9bd045c),
	.w2(32'h3a6e1e32),
	.w3(32'hb9b369c8),
	.w4(32'hb988d8bb),
	.w5(32'h3a19cbd8),
	.w6(32'hba94ded9),
	.w7(32'h393e3c08),
	.w8(32'h3a907fc0),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2881f5),
	.w1(32'h3acb260d),
	.w2(32'h3b42ef26),
	.w3(32'h3a7b2fae),
	.w4(32'h3b298c48),
	.w5(32'hba25dad5),
	.w6(32'hb9f0000f),
	.w7(32'h3b235b6f),
	.w8(32'hbaf8dde6),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38179e7d),
	.w1(32'hb994f577),
	.w2(32'h3b7b8478),
	.w3(32'hb93bed07),
	.w4(32'h3b216792),
	.w5(32'hba4a4113),
	.w6(32'hba888e27),
	.w7(32'h3acc42ec),
	.w8(32'hba9391dd),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8ff328),
	.w1(32'h3c025469),
	.w2(32'h3c25b9f1),
	.w3(32'h3a3ecdd9),
	.w4(32'h3bb57307),
	.w5(32'h3a9655e5),
	.w6(32'h3b16b70d),
	.w7(32'h3bb3372c),
	.w8(32'h388c93cf),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa1d919),
	.w1(32'hba87039f),
	.w2(32'h3b694065),
	.w3(32'hbb5788ab),
	.w4(32'h3986ea9e),
	.w5(32'hbaedb76d),
	.w6(32'hbbaf1fff),
	.w7(32'hbb1e13d8),
	.w8(32'hbaf984c4),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb02790b),
	.w1(32'hba6ea124),
	.w2(32'h3a84a298),
	.w3(32'hbb1c55b9),
	.w4(32'hb824259e),
	.w5(32'h3b474fd4),
	.w6(32'hbaa61c36),
	.w7(32'hba8af0f9),
	.w8(32'h3add1d74),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b03f8ed),
	.w1(32'h3b2579f4),
	.w2(32'h3afa3c85),
	.w3(32'h3a8fcdc1),
	.w4(32'h3a4d2c5b),
	.w5(32'hbb1b7329),
	.w6(32'h39acf3ea),
	.w7(32'h3849b203),
	.w8(32'hbadb9195),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2df936),
	.w1(32'hba9151c3),
	.w2(32'h3b5c2f95),
	.w3(32'hbad2d845),
	.w4(32'h39d62c4a),
	.w5(32'hb9e5f00e),
	.w6(32'hbb3ac635),
	.w7(32'h3a45689c),
	.w8(32'hba7419a9),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90d733d),
	.w1(32'h3a8ccfd1),
	.w2(32'h3b92e28a),
	.w3(32'h3a50ad66),
	.w4(32'h3b311107),
	.w5(32'h3abb0a60),
	.w6(32'h39cabc2e),
	.w7(32'h3a18a4d7),
	.w8(32'hba404eda),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d9f033),
	.w1(32'h3a884c25),
	.w2(32'h3bc40c93),
	.w3(32'hba8c343f),
	.w4(32'h3ba6d91b),
	.w5(32'h3ba0eb1c),
	.w6(32'hbb29b543),
	.w7(32'h3bbc8820),
	.w8(32'h3b029f74),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b0cada),
	.w1(32'hbb185703),
	.w2(32'h3b1babde),
	.w3(32'h3a97b2e3),
	.w4(32'h3b6877b7),
	.w5(32'h3a74d179),
	.w6(32'hbb251e33),
	.w7(32'h3b0f03b0),
	.w8(32'hbb160956),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad18b9e),
	.w1(32'hba042283),
	.w2(32'h3b1fa81f),
	.w3(32'h39986847),
	.w4(32'h3b190fe1),
	.w5(32'hba03d929),
	.w6(32'hbb06ced0),
	.w7(32'h3ad7b99c),
	.w8(32'hba6e6e08),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acffe72),
	.w1(32'h3a87b730),
	.w2(32'hb9f14b7d),
	.w3(32'hb8878ae6),
	.w4(32'h3917a14a),
	.w5(32'h3bcb3e80),
	.w6(32'hbb261ca2),
	.w7(32'hbaa07a6d),
	.w8(32'h3c01a995),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd2d583),
	.w1(32'h3b72f4ee),
	.w2(32'h3ae1f015),
	.w3(32'h3b38a903),
	.w4(32'h3b7707c3),
	.w5(32'h3a962e5a),
	.w6(32'h3b6645c3),
	.w7(32'h3b73b110),
	.w8(32'h3b3a57d7),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c15a879),
	.w1(32'h3c381955),
	.w2(32'h3c1e051a),
	.w3(32'h3ac347fa),
	.w4(32'h3b692dbb),
	.w5(32'h3ba9f89f),
	.w6(32'h3abec8bf),
	.w7(32'h3b20ecc2),
	.w8(32'h3b939d01),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb1722f),
	.w1(32'h3bc1b3e2),
	.w2(32'h3b891edc),
	.w3(32'h3b9952b9),
	.w4(32'h3b5bbde2),
	.w5(32'h3922ae2d),
	.w6(32'h3baa08ca),
	.w7(32'h3b05de96),
	.w8(32'h3a708847),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8bc08f),
	.w1(32'h3be8a1b3),
	.w2(32'h3c4372bc),
	.w3(32'h3c177941),
	.w4(32'h3c2c3a28),
	.w5(32'hbacc72f3),
	.w6(32'h3c23d1fb),
	.w7(32'h3c6fd3b2),
	.w8(32'hbb2abe21),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb83ca1e),
	.w1(32'hbba9f40c),
	.w2(32'hbb62c8d9),
	.w3(32'hbbc81271),
	.w4(32'hbbb98246),
	.w5(32'h3b518035),
	.w6(32'hbbd1ba73),
	.w7(32'hbb99be24),
	.w8(32'h3b23ca2f),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba480a5),
	.w1(32'h3bba85a5),
	.w2(32'h3b9e90b3),
	.w3(32'h3bf17cc9),
	.w4(32'h3bb4f98d),
	.w5(32'hbb0bc0b6),
	.w6(32'h3be7b8b0),
	.w7(32'h3bf06f59),
	.w8(32'hbb2a6832),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a9669),
	.w1(32'hba84aa21),
	.w2(32'h3ba5b1dc),
	.w3(32'hbaae6774),
	.w4(32'h3b5747a2),
	.w5(32'h3b84bea4),
	.w6(32'hbb777575),
	.w7(32'h3b2e4a11),
	.w8(32'h3b196c30),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3963c265),
	.w1(32'hbaba7154),
	.w2(32'hbb61827d),
	.w3(32'h3b2f9471),
	.w4(32'hba2e1b9f),
	.w5(32'h3b02fa4c),
	.w6(32'h3ac08913),
	.w7(32'hbac405da),
	.w8(32'h3b24c5fa),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb041f5b),
	.w1(32'hbaa7a194),
	.w2(32'hbb38b7f6),
	.w3(32'h39f8374b),
	.w4(32'hb98d05ef),
	.w5(32'h3ba15935),
	.w6(32'hbac2af1e),
	.w7(32'hba54239f),
	.w8(32'h3b36ef10),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf911be),
	.w1(32'hbadff21a),
	.w2(32'hb98d6749),
	.w3(32'h3a98e896),
	.w4(32'h3b54e1d7),
	.w5(32'hba4375fc),
	.w6(32'hb89cdc5b),
	.w7(32'h3a9005fb),
	.w8(32'hba24b385),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaea6efb),
	.w1(32'hb998b4a1),
	.w2(32'h3b1eaf01),
	.w3(32'hbaf9c1c2),
	.w4(32'h3985e714),
	.w5(32'hb9522f5f),
	.w6(32'hba94ed30),
	.w7(32'h3ac7dccb),
	.w8(32'hba96b8fa),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6b4f87),
	.w1(32'h3c7d7593),
	.w2(32'h3ca413af),
	.w3(32'h3bef18ed),
	.w4(32'h3c4a8a2d),
	.w5(32'h3b3add95),
	.w6(32'h3c0d0bf5),
	.w7(32'h3c902070),
	.w8(32'h3aeb1a6c),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae9e876),
	.w1(32'h39b0885a),
	.w2(32'h3a642aa7),
	.w3(32'h39147588),
	.w4(32'hb8b0bd61),
	.w5(32'h38d2b68c),
	.w6(32'hbb3346dd),
	.w7(32'hbb0b28dd),
	.w8(32'hb9cab8e7),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390de084),
	.w1(32'hb90d8772),
	.w2(32'h3aa38ca3),
	.w3(32'hb945f497),
	.w4(32'hb9beec02),
	.w5(32'hbad1aa02),
	.w6(32'h3b51ca38),
	.w7(32'h3a9631b9),
	.w8(32'hba3d28c0),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb349278),
	.w1(32'h3ac7ffb2),
	.w2(32'hb746310a),
	.w3(32'hbb5b7a08),
	.w4(32'hbb9ff1a9),
	.w5(32'h3b83a293),
	.w6(32'h39e63aad),
	.w7(32'h3b806e2f),
	.w8(32'h3b9f6214),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa6226e),
	.w1(32'h3ab53b93),
	.w2(32'h3b9ea4a8),
	.w3(32'hba96238e),
	.w4(32'hbb369980),
	.w5(32'h39e9f86a),
	.w6(32'hbb0e13e1),
	.w7(32'hbb781676),
	.w8(32'h3b35e532),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b08a505),
	.w1(32'hbac9869b),
	.w2(32'hbba3e89e),
	.w3(32'h3abfa44a),
	.w4(32'hbb2ba566),
	.w5(32'hbbeea9d6),
	.w6(32'h3b9a53d9),
	.w7(32'hbb8060c5),
	.w8(32'h3983afc5),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba32473b),
	.w1(32'h3a47070d),
	.w2(32'hb99778ed),
	.w3(32'hba7ce259),
	.w4(32'hbb11bef3),
	.w5(32'hbb129296),
	.w6(32'hb9a4720d),
	.w7(32'h391722ac),
	.w8(32'hbb09cfac),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab79a71),
	.w1(32'h3ab4d98b),
	.w2(32'h3b488916),
	.w3(32'hbb6e9649),
	.w4(32'h393ef1f1),
	.w5(32'h3b45c696),
	.w6(32'h3b93e6a2),
	.w7(32'h3b4c4502),
	.w8(32'h3bc909b6),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b20f41e),
	.w1(32'h3611a7a6),
	.w2(32'h3aa94410),
	.w3(32'hba323a35),
	.w4(32'hbb893adb),
	.w5(32'hbae84c74),
	.w6(32'h3b383954),
	.w7(32'hba8dbcad),
	.w8(32'hbb97f658),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8e1ce2),
	.w1(32'hb9dd4104),
	.w2(32'hbb0d7b68),
	.w3(32'hbb163503),
	.w4(32'h3a518c18),
	.w5(32'hbb1537de),
	.w6(32'h3a314dc3),
	.w7(32'hbb438c3d),
	.w8(32'hbba46381),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcdd932),
	.w1(32'hbacc7881),
	.w2(32'h3a54a429),
	.w3(32'hba85f060),
	.w4(32'hbb350b46),
	.w5(32'h3b1edc01),
	.w6(32'h3984259c),
	.w7(32'h3a0ae882),
	.w8(32'hb971e993),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af86945),
	.w1(32'h394c22db),
	.w2(32'h3a521b76),
	.w3(32'h3ad3c007),
	.w4(32'h39a01016),
	.w5(32'hbb84cdab),
	.w6(32'hbadee9f9),
	.w7(32'hbac54a06),
	.w8(32'hbb33c145),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7b8668),
	.w1(32'hba68fa65),
	.w2(32'h3b871988),
	.w3(32'h3a07842e),
	.w4(32'hbb4180fc),
	.w5(32'h3b264598),
	.w6(32'hbadbd8b1),
	.w7(32'h389c7935),
	.w8(32'hbac7bf61),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9973dd),
	.w1(32'hbb1fdca4),
	.w2(32'hbb23caa7),
	.w3(32'hbb72e24e),
	.w4(32'h3b5b17c6),
	.w5(32'h3b732d13),
	.w6(32'hbbdcea71),
	.w7(32'hbb462899),
	.w8(32'h3b23693a),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb221be4),
	.w1(32'h3a13e846),
	.w2(32'h3b41f05e),
	.w3(32'h3ae88d39),
	.w4(32'h3a017878),
	.w5(32'h3b94b8d4),
	.w6(32'h3b5dc09b),
	.w7(32'h3b0563a2),
	.w8(32'h3b83fc4f),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be5b11f),
	.w1(32'hbb468115),
	.w2(32'hbaf8c1f8),
	.w3(32'h3b6431cd),
	.w4(32'h3bb1a2e5),
	.w5(32'hbb97337b),
	.w6(32'h3ba0e46f),
	.w7(32'h3afcccbe),
	.w8(32'hbad6aaba),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb939b471),
	.w1(32'h3b33cc4c),
	.w2(32'hba1900d9),
	.w3(32'hbb745850),
	.w4(32'h3ae94404),
	.w5(32'hbb04f43f),
	.w6(32'h3b5e1c9b),
	.w7(32'h3b4c6049),
	.w8(32'hbb145632),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbc553c),
	.w1(32'hbb54c5a0),
	.w2(32'h3a10c7d2),
	.w3(32'hbb5c4962),
	.w4(32'h3ad38140),
	.w5(32'h3b942ffb),
	.w6(32'h38760744),
	.w7(32'hb99f66fc),
	.w8(32'h3b80529e),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba55e2bb),
	.w1(32'hb99ac4dd),
	.w2(32'h3b88e2e3),
	.w3(32'h3b68dbe9),
	.w4(32'h3a11d06c),
	.w5(32'h3bc657db),
	.w6(32'h3b07d336),
	.w7(32'h39bdd17b),
	.w8(32'h3b1b22ab),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b10a6b5),
	.w1(32'h3bec54ae),
	.w2(32'h3bb69a43),
	.w3(32'h3bc00a0a),
	.w4(32'h3bec012f),
	.w5(32'hbb0b1b3f),
	.w6(32'h3b358a61),
	.w7(32'h3b9993c4),
	.w8(32'hb95b8a36),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb62a7a3),
	.w1(32'hbb04970b),
	.w2(32'h3aa5bdb8),
	.w3(32'hb9431429),
	.w4(32'hbb1c8aff),
	.w5(32'h3b2bf4df),
	.w6(32'h3b073646),
	.w7(32'hba6f7db1),
	.w8(32'h39ec4088),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3920f907),
	.w1(32'hbb135494),
	.w2(32'hb9ef5215),
	.w3(32'h38e805f1),
	.w4(32'h3b03cb8a),
	.w5(32'hbacddf57),
	.w6(32'hbaf2ff6c),
	.w7(32'hb9a50199),
	.w8(32'hbb0fa2fc),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1b1964),
	.w1(32'hba5a65e5),
	.w2(32'h3a9912c1),
	.w3(32'hba209bc0),
	.w4(32'h3adbe34f),
	.w5(32'h3ad0ed14),
	.w6(32'hbbe7a1c4),
	.w7(32'hbb567bca),
	.w8(32'h3acdbab4),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h380aecec),
	.w1(32'hbac4d4c8),
	.w2(32'hba87e44f),
	.w3(32'hba837e34),
	.w4(32'h3a38fc1b),
	.w5(32'h3a967644),
	.w6(32'h3aa661f1),
	.w7(32'h3a8c89b1),
	.w8(32'h3b112cf8),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0f83eb),
	.w1(32'hbbff0097),
	.w2(32'hba56f028),
	.w3(32'h3b0b5938),
	.w4(32'h3ac64530),
	.w5(32'hbadfe91e),
	.w6(32'h3a644f17),
	.w7(32'h3b1825d8),
	.w8(32'h3bc1c359),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97e9721),
	.w1(32'hbac3a978),
	.w2(32'hbab92969),
	.w3(32'hbb230e0b),
	.w4(32'hbbad82af),
	.w5(32'hbba3e46f),
	.w6(32'h3aa42466),
	.w7(32'hbbba763b),
	.w8(32'hbb5a811b),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6793b5),
	.w1(32'hbb39e957),
	.w2(32'hbb7f90cf),
	.w3(32'h3b0cbdec),
	.w4(32'h3a7d6e61),
	.w5(32'hb9480c8a),
	.w6(32'h3a701e94),
	.w7(32'h3a93b73c),
	.w8(32'h3b1c22bb),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b195eee),
	.w1(32'h3b4b9271),
	.w2(32'hb95b162f),
	.w3(32'hb89e6a14),
	.w4(32'hbac2eebb),
	.w5(32'hbb2c23d2),
	.w6(32'hbad8d957),
	.w7(32'hbbe078cb),
	.w8(32'hbb56d194),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaea5000),
	.w1(32'h3910b391),
	.w2(32'h3aa2aacb),
	.w3(32'h3a6bf01e),
	.w4(32'h3a9a16c5),
	.w5(32'hbb8983b7),
	.w6(32'h3a09cbc2),
	.w7(32'h3ae98f93),
	.w8(32'hbb5f6bf6),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9da217),
	.w1(32'h3a938f16),
	.w2(32'h3b75729f),
	.w3(32'h398b7a47),
	.w4(32'hbb076f52),
	.w5(32'h3971939b),
	.w6(32'h3b5a4f74),
	.w7(32'h3b230838),
	.w8(32'hba0fa941),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb44a91b),
	.w1(32'h3ae41288),
	.w2(32'hbb6cb003),
	.w3(32'hb9383dcd),
	.w4(32'hbb204f93),
	.w5(32'h3c02ef64),
	.w6(32'h3b329d0a),
	.w7(32'hb9ba07dc),
	.w8(32'h3c8991aa),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c38c6ef),
	.w1(32'h3a932405),
	.w2(32'h3b458cb5),
	.w3(32'h3c5ce52c),
	.w4(32'h3bc43ec3),
	.w5(32'hb9792b80),
	.w6(32'h3c77b7f3),
	.w7(32'h3b20044e),
	.w8(32'h3b5a8186),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf7b124),
	.w1(32'h3acff70c),
	.w2(32'h39ba4c11),
	.w3(32'h3b850c6f),
	.w4(32'h39d21bfd),
	.w5(32'h3ae13280),
	.w6(32'h3c117650),
	.w7(32'h3a73c869),
	.w8(32'hbb046589),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396c7942),
	.w1(32'hbab56195),
	.w2(32'hb94c13b3),
	.w3(32'hbb216a28),
	.w4(32'h3ab39e2c),
	.w5(32'h3ae6192d),
	.w6(32'hba904563),
	.w7(32'h398e8322),
	.w8(32'h3b80961c),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8b621b),
	.w1(32'h3abae4f1),
	.w2(32'h3af5560b),
	.w3(32'h3b05ad24),
	.w4(32'h3ab09915),
	.w5(32'hbb189351),
	.w6(32'h3a7e44e7),
	.w7(32'hba5bf122),
	.w8(32'hba353efb),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4879a4),
	.w1(32'hbb8be18b),
	.w2(32'hbbc36b42),
	.w3(32'hbb2e4494),
	.w4(32'hbba9651d),
	.w5(32'hba1a788d),
	.w6(32'hbb97faf3),
	.w7(32'hbc1bf442),
	.w8(32'hb8c9e928),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb16e453),
	.w1(32'h3a9d3aec),
	.w2(32'h3b410115),
	.w3(32'h39143688),
	.w4(32'hbb5453d4),
	.w5(32'h3b8e6f7f),
	.w6(32'hb850eb5c),
	.w7(32'hb99d7c8a),
	.w8(32'h3ab653f8),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba564698),
	.w1(32'h3b149fad),
	.w2(32'h3b845b1c),
	.w3(32'h39b79e6f),
	.w4(32'hbb0da44c),
	.w5(32'h3c7852df),
	.w6(32'h3b8254e6),
	.w7(32'h3b37e2ce),
	.w8(32'h3c6e1412),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc6895c),
	.w1(32'hbc1734fe),
	.w2(32'hbb50a1d7),
	.w3(32'h3c2e16e8),
	.w4(32'h3be70c4e),
	.w5(32'h3be65413),
	.w6(32'hbbd0c6d5),
	.w7(32'hbbe74268),
	.w8(32'h3b89cd74),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9464c6),
	.w1(32'h3b45200a),
	.w2(32'h3b801017),
	.w3(32'h3bc67ff8),
	.w4(32'h3bcbf7a8),
	.w5(32'hbb4d266a),
	.w6(32'h3b8d459e),
	.w7(32'h3b39bfce),
	.w8(32'hb981675a),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb015c49),
	.w1(32'h393712ee),
	.w2(32'h3b155541),
	.w3(32'h3b325388),
	.w4(32'hbb8e06e1),
	.w5(32'hbaa9a0f5),
	.w6(32'h3ae03382),
	.w7(32'hb9cb4d8d),
	.w8(32'h3b44a2a1),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0615a1),
	.w1(32'hbb121b16),
	.w2(32'hb8093d3c),
	.w3(32'hba4f99dc),
	.w4(32'hbb685fc7),
	.w5(32'h3b3d606f),
	.w6(32'h3a4c63f3),
	.w7(32'hbb2c6353),
	.w8(32'hbacd36c8),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bacea12),
	.w1(32'h3b661b00),
	.w2(32'hbaf1aac3),
	.w3(32'hbb6df3b5),
	.w4(32'hbb0f711d),
	.w5(32'hbbf9450e),
	.w6(32'h39612609),
	.w7(32'h3b4da04c),
	.w8(32'hba9f9796),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8d5ef7),
	.w1(32'hbbddd2a3),
	.w2(32'hbba4ea09),
	.w3(32'h36d075f8),
	.w4(32'hbb98f1b3),
	.w5(32'hbba6a191),
	.w6(32'hbb365a6b),
	.w7(32'hbc1b417d),
	.w8(32'hbb01ef6f),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb989a46),
	.w1(32'h39021474),
	.w2(32'h398a2fc7),
	.w3(32'h3aa2195f),
	.w4(32'h3b4eb636),
	.w5(32'h3bb2851a),
	.w6(32'h3aafd31a),
	.w7(32'h3a694a82),
	.w8(32'h3b044ec4),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3bf97b),
	.w1(32'hb9c544a1),
	.w2(32'hbad7d2af),
	.w3(32'hbab2c04f),
	.w4(32'h3b0e9182),
	.w5(32'hba2149c4),
	.w6(32'hbb827af4),
	.w7(32'hba1bf5cb),
	.w8(32'h3ad8a12d),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a780792),
	.w1(32'hbb28845d),
	.w2(32'hb908cf78),
	.w3(32'h3a48e56b),
	.w4(32'hbade42d1),
	.w5(32'h3b07d6ae),
	.w6(32'h3b62ae9a),
	.w7(32'h3b4e8fbc),
	.w8(32'hbb106b2f),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2e069f),
	.w1(32'h3bbb2fd1),
	.w2(32'h3a0ee36a),
	.w3(32'h3b39ff49),
	.w4(32'hbb32a0ff),
	.w5(32'hb70ecd6b),
	.w6(32'h3c0d166a),
	.w7(32'h3b857dfb),
	.w8(32'hb91b570c),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afd18aa),
	.w1(32'h3a1f8bdc),
	.w2(32'hba28b93f),
	.w3(32'h3a2bb365),
	.w4(32'hb993e471),
	.w5(32'h3890727e),
	.w6(32'h3b045545),
	.w7(32'h396d771b),
	.w8(32'hba5c1973),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d7a918),
	.w1(32'hba7cf3c4),
	.w2(32'hbafb46b7),
	.w3(32'hbace1810),
	.w4(32'hba95edc9),
	.w5(32'hbb88252e),
	.w6(32'hb872bba8),
	.w7(32'h3a5a9e6d),
	.w8(32'hbb865a61),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6d59b7),
	.w1(32'h3ae677d6),
	.w2(32'h3b98ae87),
	.w3(32'hb8611bdc),
	.w4(32'h3ae7e5a1),
	.w5(32'hb6536247),
	.w6(32'h3b194417),
	.w7(32'h3b0f4f79),
	.w8(32'hb91938ac),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb030871),
	.w1(32'hbb9ee333),
	.w2(32'h3b198ec1),
	.w3(32'h3a310c80),
	.w4(32'h3b42c5a0),
	.w5(32'h3b22d437),
	.w6(32'h39ca1afa),
	.w7(32'h3bcf39ff),
	.w8(32'h3affba62),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b45615d),
	.w1(32'h3c0d434d),
	.w2(32'h3c04d166),
	.w3(32'h3b381c07),
	.w4(32'h3bc73bc1),
	.w5(32'hbb89d262),
	.w6(32'h3b3863f1),
	.w7(32'h3ba0d5f9),
	.w8(32'hba6e2610),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abe580d),
	.w1(32'hb80fe595),
	.w2(32'hbb3d6ff8),
	.w3(32'hbbd1de6a),
	.w4(32'hba75a018),
	.w5(32'h3b6c88d6),
	.w6(32'h3aad05fe),
	.w7(32'hb97c9649),
	.w8(32'h3bb9afe9),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb95db34),
	.w1(32'hbc110216),
	.w2(32'hbb4f987d),
	.w3(32'h3ba2239c),
	.w4(32'hbb85390b),
	.w5(32'h3b58b689),
	.w6(32'hba3f7208),
	.w7(32'hbbc44dcb),
	.w8(32'h3b3a7538),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb19d82d),
	.w1(32'hb91ee174),
	.w2(32'h3ba479c9),
	.w3(32'hbb82b68e),
	.w4(32'hbb2872dd),
	.w5(32'h3b24d928),
	.w6(32'hbb4bf06e),
	.w7(32'hbadd84d7),
	.w8(32'hbb7a8543),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb03391c),
	.w1(32'h3af7f922),
	.w2(32'hba722027),
	.w3(32'hba64013d),
	.w4(32'hbab9772c),
	.w5(32'h3b0a22ba),
	.w6(32'hbb0370dd),
	.w7(32'h3a60f3cd),
	.w8(32'h39121892),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab8b66e),
	.w1(32'h3abef1c9),
	.w2(32'h3989e74c),
	.w3(32'hba57eea5),
	.w4(32'hb8bb38fc),
	.w5(32'h3a9c61a1),
	.w6(32'hba9d2b25),
	.w7(32'h3a025a1c),
	.w8(32'h3b5830f6),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b66cd2c),
	.w1(32'h3b665445),
	.w2(32'h3bc93f9b),
	.w3(32'h3c0b199d),
	.w4(32'h3b955810),
	.w5(32'hbb947b3d),
	.w6(32'h3c05eaa0),
	.w7(32'h3bcff42b),
	.w8(32'hbac6c682),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a658710),
	.w1(32'h3b67e0ef),
	.w2(32'h3b0d0900),
	.w3(32'h3a01e33c),
	.w4(32'hbac34e5f),
	.w5(32'hba28d86f),
	.w6(32'h3b731da5),
	.w7(32'h3b057f4b),
	.w8(32'hbacba201),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1e7c26),
	.w1(32'hbbe857e7),
	.w2(32'hba903ae0),
	.w3(32'h3ae2d609),
	.w4(32'h39883d44),
	.w5(32'hba117a46),
	.w6(32'hbb111f13),
	.w7(32'h39dce576),
	.w8(32'h3b9b7c31),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb545358),
	.w1(32'hbb6cf4e2),
	.w2(32'hbae59f41),
	.w3(32'hbb1ea4fb),
	.w4(32'hbba75de5),
	.w5(32'hbbd0e519),
	.w6(32'hbc329c2d),
	.w7(32'hbbb76fbc),
	.w8(32'hbc07046a),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2b02c9),
	.w1(32'h3b1e9a7f),
	.w2(32'hbb0ad007),
	.w3(32'hbb232f08),
	.w4(32'h38b3f340),
	.w5(32'h3a88403d),
	.w6(32'h3a0c935e),
	.w7(32'hbacdb160),
	.w8(32'h3b8dc948),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb124945),
	.w1(32'h3b766914),
	.w2(32'hba07ca64),
	.w3(32'h3adf6dd3),
	.w4(32'hbb0c4a87),
	.w5(32'hba06170a),
	.w6(32'h3aba5b39),
	.w7(32'h392bdba2),
	.w8(32'hb8e55b21),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba56cf52),
	.w1(32'h39abfa07),
	.w2(32'hba1e8696),
	.w3(32'h3b1e3a58),
	.w4(32'hbb0a10e4),
	.w5(32'hbb8fef80),
	.w6(32'h3b6af402),
	.w7(32'hb9db7963),
	.w8(32'hbb31f5d5),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba678783),
	.w1(32'h3a8efffd),
	.w2(32'h3b260d66),
	.w3(32'hbb66a8a6),
	.w4(32'hbb89b666),
	.w5(32'h3a8e8b2d),
	.w6(32'hba064155),
	.w7(32'hb98b8beb),
	.w8(32'hba2a5403),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2f65b4),
	.w1(32'hbb8b5fca),
	.w2(32'hbb83a602),
	.w3(32'hbb383bc6),
	.w4(32'hbb4254c4),
	.w5(32'hbb2333b0),
	.w6(32'h38e3388a),
	.w7(32'hbb1e20de),
	.w8(32'h3a2012dc),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb997a83),
	.w1(32'hbac92114),
	.w2(32'hbaf361e1),
	.w3(32'hbba5f836),
	.w4(32'hbbb4458c),
	.w5(32'h3a67f6a8),
	.w6(32'hbb4f0a26),
	.w7(32'hbae3509c),
	.w8(32'h3a44cf97),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3c56d7),
	.w1(32'h3b3957e9),
	.w2(32'h3b58ae0f),
	.w3(32'hbb50468a),
	.w4(32'hbbba8809),
	.w5(32'hbaa33360),
	.w6(32'hba01eacd),
	.w7(32'h3ac39b6c),
	.w8(32'h3b8c2986),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa1f0c0),
	.w1(32'h3a7d89f8),
	.w2(32'h3a0adf1d),
	.w3(32'hba69ba30),
	.w4(32'hbb12e592),
	.w5(32'h3aeb9eda),
	.w6(32'h3b52c5bd),
	.w7(32'hbb7bde7a),
	.w8(32'h3b821b58),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b70e64a),
	.w1(32'h3b5554c2),
	.w2(32'h3bc3027d),
	.w3(32'h3b470ae1),
	.w4(32'h3b7df160),
	.w5(32'hbbab66cd),
	.w6(32'h3bf5c733),
	.w7(32'h3bea20db),
	.w8(32'hb9dd8de7),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5b76b0),
	.w1(32'h3b4d7f05),
	.w2(32'hbb572eb2),
	.w3(32'h3aaba612),
	.w4(32'h3aee5725),
	.w5(32'hbaf8fa53),
	.w6(32'h3bd429c2),
	.w7(32'h3b58d526),
	.w8(32'hbac10578),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb896847),
	.w1(32'h3a2e0b24),
	.w2(32'h3aadb3dd),
	.w3(32'hbb0a6c7b),
	.w4(32'hbad2d35a),
	.w5(32'hbbafe1e1),
	.w6(32'hbb384eed),
	.w7(32'h3a24ca6c),
	.w8(32'hbb3b0ce1),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf6c923),
	.w1(32'hbb711e3f),
	.w2(32'hb9867ca3),
	.w3(32'hbc056341),
	.w4(32'hbb677990),
	.w5(32'hba3b2b9b),
	.w6(32'hbbfb5f3d),
	.w7(32'hbb9e0fab),
	.w8(32'hbac1f398),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bc97c1),
	.w1(32'h3a712be7),
	.w2(32'h3a05c200),
	.w3(32'hbb5be206),
	.w4(32'hba0874fc),
	.w5(32'hbb6be52c),
	.w6(32'h3a8ee00e),
	.w7(32'hb94dd4c1),
	.w8(32'hbab90687),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb93a46a),
	.w1(32'hbb3b40ca),
	.w2(32'h3b1a38e5),
	.w3(32'hbbcdfafe),
	.w4(32'hbb861827),
	.w5(32'h39e58037),
	.w6(32'hbbb5e58a),
	.w7(32'hbaf3e946),
	.w8(32'hbb49bb6d),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b924f),
	.w1(32'h397f9700),
	.w2(32'h3bdfc9b3),
	.w3(32'hbb872962),
	.w4(32'hbb881d6d),
	.w5(32'hba1f0459),
	.w6(32'h38b42a8b),
	.w7(32'h3b12e25c),
	.w8(32'hbb0441a1),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba682e6b),
	.w1(32'h3ae38fdc),
	.w2(32'h3b36aa52),
	.w3(32'hbb3557a6),
	.w4(32'hbab66136),
	.w5(32'h3bda6771),
	.w6(32'hbaadebcf),
	.w7(32'hba055d37),
	.w8(32'h3bca1a5d),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9421b0),
	.w1(32'h3bc2e6e5),
	.w2(32'h3b631349),
	.w3(32'h3baa02bc),
	.w4(32'h3bd67472),
	.w5(32'hba63f47b),
	.w6(32'h3b553918),
	.w7(32'h3b685d6a),
	.w8(32'h3b5fb494),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bbd583),
	.w1(32'hbb5d39a1),
	.w2(32'hba9c5f9b),
	.w3(32'h3b312350),
	.w4(32'hbad92624),
	.w5(32'h3b8da054),
	.w6(32'hbb5fddd3),
	.w7(32'hbbb89894),
	.w8(32'h3b456e90),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba39d78),
	.w1(32'h3be18b1d),
	.w2(32'h3ba611de),
	.w3(32'h3aeb2be8),
	.w4(32'h3bbfc256),
	.w5(32'h3bc198cc),
	.w6(32'hb8dcbf04),
	.w7(32'h3b72c3b9),
	.w8(32'h3b7210bd),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3993eec0),
	.w1(32'h3b534d0c),
	.w2(32'h3b16a769),
	.w3(32'h3b12372c),
	.w4(32'h3aed94a2),
	.w5(32'h3a6bc68d),
	.w6(32'h3b2c23fd),
	.w7(32'h3aadb260),
	.w8(32'h39af7e11),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb73d0f08),
	.w1(32'h3b168150),
	.w2(32'h3adea697),
	.w3(32'hb8ffecf4),
	.w4(32'h3a1ed902),
	.w5(32'hba9cd719),
	.w6(32'h3b180dbe),
	.w7(32'h3ad02dba),
	.w8(32'hb974f9ac),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ed5d70),
	.w1(32'hbbc4eca1),
	.w2(32'hbb46ae7d),
	.w3(32'hbbcdd0bc),
	.w4(32'hbb531a98),
	.w5(32'h3a906c42),
	.w6(32'hba47fcbc),
	.w7(32'hbb45b037),
	.w8(32'hbb47bec8),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb37193d),
	.w1(32'hbb8a9b74),
	.w2(32'h3b229b34),
	.w3(32'hbb8eeb5a),
	.w4(32'hb9918024),
	.w5(32'hbb524e75),
	.w6(32'hbb0c2150),
	.w7(32'h3b919314),
	.w8(32'hbb41e8da),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad03220),
	.w1(32'h3b3d68db),
	.w2(32'h3ae7c655),
	.w3(32'hba73c622),
	.w4(32'hba3c77e7),
	.w5(32'hbb3b43f9),
	.w6(32'h3b480865),
	.w7(32'h3acc81ae),
	.w8(32'hba3f5185),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0cef07),
	.w1(32'h3b63d20b),
	.w2(32'h3b52bfd8),
	.w3(32'hb6baf264),
	.w4(32'hbb2d8e4d),
	.w5(32'hbb023ef2),
	.w6(32'h3abfd0bc),
	.w7(32'h39d673eb),
	.w8(32'hbac963f8),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7f20ed),
	.w1(32'h3b59c1c1),
	.w2(32'hb91ad311),
	.w3(32'h3b721fa2),
	.w4(32'h3adf5659),
	.w5(32'hbbd1d6d3),
	.w6(32'h3b0a0eb4),
	.w7(32'h3ade01f6),
	.w8(32'hba878f00),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b091b1a),
	.w1(32'hbb4c2bca),
	.w2(32'h3b30659b),
	.w3(32'hbb56e72b),
	.w4(32'h3a262eb5),
	.w5(32'h3bc9a4bf),
	.w6(32'h3ab673f0),
	.w7(32'h3b4dc1c2),
	.w8(32'h3a51dcb9),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8ee449),
	.w1(32'h3bbc0ccd),
	.w2(32'h3b8503be),
	.w3(32'h3b3c6bf9),
	.w4(32'h3bc5fd29),
	.w5(32'hbb2e1a42),
	.w6(32'hb9bfbdf2),
	.w7(32'h3ba394cd),
	.w8(32'hbb7cec8e),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac28138),
	.w1(32'h3c160234),
	.w2(32'h3bf7d452),
	.w3(32'hbc12e33d),
	.w4(32'hbbe00192),
	.w5(32'h39cde9aa),
	.w6(32'hbba1ef91),
	.w7(32'hbbc9cc5c),
	.w8(32'h3ba21772),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1bebce),
	.w1(32'hba8e0951),
	.w2(32'hbaf4e527),
	.w3(32'hbb3ae553),
	.w4(32'h3b62ed03),
	.w5(32'hbbab6789),
	.w6(32'hb9000d1b),
	.w7(32'h3a5d9d6c),
	.w8(32'hbb8a5d11),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba75ed52),
	.w1(32'h3aa7c257),
	.w2(32'h3ae4baae),
	.w3(32'hba9f8dd3),
	.w4(32'hbb0b246a),
	.w5(32'hbb2938d2),
	.w6(32'h3a8a1204),
	.w7(32'h3a1654f1),
	.w8(32'h3aaa332f),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa1b94e),
	.w1(32'h39327298),
	.w2(32'hb9f8eada),
	.w3(32'hba7208b6),
	.w4(32'hbb293e70),
	.w5(32'hbb4f5957),
	.w6(32'h3b44ee1d),
	.w7(32'h3a87c703),
	.w8(32'hbaa92334),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9928288),
	.w1(32'hba130f37),
	.w2(32'hbb1d65d8),
	.w3(32'h3a88f6cf),
	.w4(32'hbb1631c3),
	.w5(32'hbb5d81ac),
	.w6(32'h3a58a9c9),
	.w7(32'hbb1d2038),
	.w8(32'hbb95a83d),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3ebf42),
	.w1(32'h3ada10bd),
	.w2(32'h3a0a3dff),
	.w3(32'h3b6186fb),
	.w4(32'h3932fca0),
	.w5(32'hbb80c28a),
	.w6(32'h3b22e3ab),
	.w7(32'h3ab45bdd),
	.w8(32'h39603ce6),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6f195f),
	.w1(32'h3a5f53be),
	.w2(32'hbab889ea),
	.w3(32'hbb3d4c1a),
	.w4(32'hbba5d465),
	.w5(32'h3bc79b17),
	.w6(32'h3b9216d0),
	.w7(32'hba1b7519),
	.w8(32'h3bdaf635),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2aa2b9),
	.w1(32'hbbc92ee7),
	.w2(32'hba9c51d0),
	.w3(32'hba1e8f1d),
	.w4(32'h3aacd874),
	.w5(32'hbab40877),
	.w6(32'hbabd82f4),
	.w7(32'hbb20220a),
	.w8(32'hbb569ad8),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe12ace),
	.w1(32'hbc05c538),
	.w2(32'hbbb7be38),
	.w3(32'hbba67a31),
	.w4(32'hbb52dc7b),
	.w5(32'h3b04a8e1),
	.w6(32'hbc744e2c),
	.w7(32'hbc0cd568),
	.w8(32'h3a049574),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb1f073),
	.w1(32'hbb0d2353),
	.w2(32'hbb1d9f12),
	.w3(32'h3b62d193),
	.w4(32'hba598b68),
	.w5(32'h3af4e981),
	.w6(32'h3629e96a),
	.w7(32'hba52d2e6),
	.w8(32'hb99ccbf7),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2dfc19),
	.w1(32'hb9bf0b20),
	.w2(32'h3b1eb3a6),
	.w3(32'hb97f21fa),
	.w4(32'hbb056715),
	.w5(32'hba405a61),
	.w6(32'hbb05bc98),
	.w7(32'hbaf99f42),
	.w8(32'h39b5eda1),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba880b47),
	.w1(32'hbad44ddb),
	.w2(32'hbaa23ed9),
	.w3(32'hbb1269cd),
	.w4(32'hbb344e4f),
	.w5(32'h3be1e727),
	.w6(32'hbb10ac4c),
	.w7(32'hbb277184),
	.w8(32'h3b9a7066),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0acb16),
	.w1(32'hbc14c767),
	.w2(32'hba9016c1),
	.w3(32'h3ba0eae4),
	.w4(32'hba337d54),
	.w5(32'h3b525d8f),
	.w6(32'h3b892715),
	.w7(32'hbaf57c98),
	.w8(32'h3b5327d6),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac17451),
	.w1(32'hba7e3a9a),
	.w2(32'hbb5e2f77),
	.w3(32'h3abce84a),
	.w4(32'h3ac7770f),
	.w5(32'hbb7ecbe7),
	.w6(32'h3b2f8664),
	.w7(32'hbbb396e5),
	.w8(32'hbad5e115),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac8083f),
	.w1(32'hb866aa14),
	.w2(32'h37eaf406),
	.w3(32'hb991193f),
	.w4(32'hb99768a1),
	.w5(32'hba94557f),
	.w6(32'hba2abab3),
	.w7(32'h37e69d36),
	.w8(32'h3b151fe9),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfbac05),
	.w1(32'hbb7e6a14),
	.w2(32'hbb4f44f8),
	.w3(32'hbb8d8297),
	.w4(32'hbb5d7805),
	.w5(32'hbbd3e8e7),
	.w6(32'h3b973bdc),
	.w7(32'h3a854e23),
	.w8(32'hbb3d238a),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab786b5),
	.w1(32'hbb511d35),
	.w2(32'hbbbae8cb),
	.w3(32'hbabc0ad8),
	.w4(32'hbb5ef157),
	.w5(32'hbb3f3605),
	.w6(32'hbad438fd),
	.w7(32'hbbb904fc),
	.w8(32'h3b0c530b),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3c9c91),
	.w1(32'hbaac9548),
	.w2(32'hbb57f00c),
	.w3(32'hb9b723cd),
	.w4(32'h3a9e6f5d),
	.w5(32'h39325e98),
	.w6(32'h3b6be478),
	.w7(32'hba6c7ffb),
	.w8(32'h3a255891),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b7ff56),
	.w1(32'hbaafc2e5),
	.w2(32'hbad34fd2),
	.w3(32'hba800566),
	.w4(32'hbaa62768),
	.w5(32'h3b26ae6f),
	.w6(32'h3a8b0ad8),
	.w7(32'hb92e1d97),
	.w8(32'h3bf4d9c7),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be42eb6),
	.w1(32'hba0f9c5e),
	.w2(32'h36651de9),
	.w3(32'h3b944075),
	.w4(32'h3b706e79),
	.w5(32'h3af0ed7a),
	.w6(32'h3b007872),
	.w7(32'hbb14bf33),
	.w8(32'h3ac105fe),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7297844),
	.w1(32'hbaf1048e),
	.w2(32'h3ab99acc),
	.w3(32'h3b0b2826),
	.w4(32'hbb6c6bd0),
	.w5(32'h3bf47a97),
	.w6(32'h3b404e38),
	.w7(32'hbafad2da),
	.w8(32'h3ba18a43),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b05a0f4),
	.w1(32'hbb8048f2),
	.w2(32'h3b2dd023),
	.w3(32'h3c010206),
	.w4(32'h3c16e1b3),
	.w5(32'h3b3c45c8),
	.w6(32'hbc02aecf),
	.w7(32'hbb332850),
	.w8(32'h3b94c8e2),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39aa8b91),
	.w1(32'h3a84fa55),
	.w2(32'h39cf6a10),
	.w3(32'h3ae5dde1),
	.w4(32'h37730f3a),
	.w5(32'h3a007f39),
	.w6(32'h391d23ac),
	.w7(32'hba43cccc),
	.w8(32'h3a74cae3),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba21d869),
	.w1(32'hbac6ea9c),
	.w2(32'hbac14815),
	.w3(32'h3ae116df),
	.w4(32'h3a98f9fc),
	.w5(32'hbb83e82e),
	.w6(32'h3b81915f),
	.w7(32'hbad8714a),
	.w8(32'h3a26af69),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a448f7a),
	.w1(32'hba9d38c4),
	.w2(32'hbb45b764),
	.w3(32'h3b121fac),
	.w4(32'hbab7793d),
	.w5(32'hbaab817b),
	.w6(32'h3af9d2c6),
	.w7(32'h3a9070a6),
	.w8(32'h3a353d4a),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b00071a),
	.w1(32'h3af0fe57),
	.w2(32'hba1a6eef),
	.w3(32'hbb0ce2eb),
	.w4(32'hb9d6279b),
	.w5(32'hbb9de059),
	.w6(32'h3b6058d3),
	.w7(32'h3ab43ac2),
	.w8(32'h3ae31623),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb68945f),
	.w1(32'hbb7fddbf),
	.w2(32'h3acb3787),
	.w3(32'hba9c9b6a),
	.w4(32'h3983fcc9),
	.w5(32'h3bb556f5),
	.w6(32'hbb1c73dd),
	.w7(32'hbbcfbbde),
	.w8(32'hb7a4d4b1),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e16c68),
	.w1(32'hbaf29c6b),
	.w2(32'hbb36d3c3),
	.w3(32'hbb5972a1),
	.w4(32'hbb1889fd),
	.w5(32'hbb428c66),
	.w6(32'hbb550361),
	.w7(32'h3adc672b),
	.w8(32'hb9dc3038),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7d234c),
	.w1(32'hbb2bb7d7),
	.w2(32'hbb874aa0),
	.w3(32'h3ab7d467),
	.w4(32'h3a5ff063),
	.w5(32'h3b074233),
	.w6(32'h399ef60a),
	.w7(32'hbb09c079),
	.w8(32'hbaabc127),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb956e87e),
	.w1(32'h3b8290ce),
	.w2(32'h3b19d8c3),
	.w3(32'hba269653),
	.w4(32'hba05f640),
	.w5(32'h3ae4cb1f),
	.w6(32'h3b09167e),
	.w7(32'h3b139afc),
	.w8(32'h3ab4cac7),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5047c3),
	.w1(32'hbc29716c),
	.w2(32'hb9a5482a),
	.w3(32'h3c28a624),
	.w4(32'hba80fdde),
	.w5(32'h3ac123ac),
	.w6(32'h3b402921),
	.w7(32'hb9597c4c),
	.w8(32'h3b2885fc),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf34cb1),
	.w1(32'hba13857f),
	.w2(32'h3b91f02d),
	.w3(32'h3b40fe87),
	.w4(32'h384371d6),
	.w5(32'h39c07e90),
	.w6(32'h3b896af7),
	.w7(32'h3b2e767e),
	.w8(32'h3ad34777),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1e7aa6),
	.w1(32'hba1b6d23),
	.w2(32'hba3b6c30),
	.w3(32'h3b8ebf87),
	.w4(32'hbb268700),
	.w5(32'hbb90e959),
	.w6(32'h3b3bbaaf),
	.w7(32'hba99363d),
	.w8(32'hbb393241),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b0160),
	.w1(32'hba718d41),
	.w2(32'hbb89e9e9),
	.w3(32'hbb96b8c6),
	.w4(32'hbb1e1f99),
	.w5(32'hb9877a66),
	.w6(32'hbb6d69c6),
	.w7(32'hba1f3f04),
	.w8(32'hbaa5b512),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3dc896),
	.w1(32'hba9143b9),
	.w2(32'h3b1c6ba7),
	.w3(32'hbb2d6a59),
	.w4(32'h3af1fea9),
	.w5(32'h396cb93a),
	.w6(32'hbb179f60),
	.w7(32'h3b23642c),
	.w8(32'h3b16a6d3),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa1844d),
	.w1(32'hbb039003),
	.w2(32'h3a35af58),
	.w3(32'h3a6e6d40),
	.w4(32'hbb95d3a5),
	.w5(32'h391ad204),
	.w6(32'hb920f0d2),
	.w7(32'h376b3eb7),
	.w8(32'hbbb069d5),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa8be0a),
	.w1(32'hbb1280c6),
	.w2(32'hbaf18f9f),
	.w3(32'hbba5bebe),
	.w4(32'hba80ea18),
	.w5(32'hbb6c41a3),
	.w6(32'hbb34e04b),
	.w7(32'h3ae8aa5e),
	.w8(32'h3a819e4b),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa756a4),
	.w1(32'h3b9935bb),
	.w2(32'h3ae6a433),
	.w3(32'h3b8fecb2),
	.w4(32'h3bc43474),
	.w5(32'hbb69b643),
	.w6(32'h3bad90b7),
	.w7(32'h3b7019e4),
	.w8(32'h3a95e810),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc8280a),
	.w1(32'h3b8f1d1f),
	.w2(32'hbb7ad1de),
	.w3(32'h3b034436),
	.w4(32'hbaf2500a),
	.w5(32'hba9d72f9),
	.w6(32'h3b0f4615),
	.w7(32'hb96fddc5),
	.w8(32'hba28f396),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb939078b),
	.w1(32'hb9253b83),
	.w2(32'hba445e93),
	.w3(32'h3901c171),
	.w4(32'hb95a7ed7),
	.w5(32'hba521050),
	.w6(32'hb99d0fef),
	.w7(32'hb9460fef),
	.w8(32'hba65dbda),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a820a4b),
	.w1(32'hb8bcf935),
	.w2(32'hb8dadc54),
	.w3(32'hb9804df4),
	.w4(32'h3a729a23),
	.w5(32'h3ac0f3a2),
	.w6(32'hb9e87e3b),
	.w7(32'h3a8f363e),
	.w8(32'h3b6d7aff),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aca951f),
	.w1(32'h3a8f7e27),
	.w2(32'h3ad8ac2d),
	.w3(32'h3afae71e),
	.w4(32'h39f8a29e),
	.w5(32'hbb56403d),
	.w6(32'h3b9d586e),
	.w7(32'h3b6117fa),
	.w8(32'hbaecdfa7),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba037a61),
	.w1(32'hb9146ed4),
	.w2(32'h3aaa2bf9),
	.w3(32'hbacbc485),
	.w4(32'h3b0531e5),
	.w5(32'hba595bb4),
	.w6(32'hba26b36c),
	.w7(32'h3a6b76ce),
	.w8(32'hba3fc713),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a35619a),
	.w1(32'h3979a268),
	.w2(32'hb988eec7),
	.w3(32'h3b62be52),
	.w4(32'hbb20d112),
	.w5(32'hbb10034c),
	.w6(32'h3b846c2c),
	.w7(32'h37177789),
	.w8(32'hbb2fb8c6),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaed8687),
	.w1(32'hbb9844ca),
	.w2(32'hbb21d933),
	.w3(32'hbb97a92a),
	.w4(32'hbb08ffbb),
	.w5(32'h3b244742),
	.w6(32'hbbef4f8d),
	.w7(32'hbb8aacad),
	.w8(32'h3b54394a),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba13d75a),
	.w1(32'hbb02fb3e),
	.w2(32'hba32dc48),
	.w3(32'h3ac3b345),
	.w4(32'hba0c19d6),
	.w5(32'h39d095be),
	.w6(32'h3aaa6802),
	.w7(32'hbab7d82a),
	.w8(32'hba71a919),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bef4a4),
	.w1(32'hba3f2fb5),
	.w2(32'h3a23cd8b),
	.w3(32'hba4564e6),
	.w4(32'hb9a6960a),
	.w5(32'h3a9aef00),
	.w6(32'hba07f182),
	.w7(32'hb9f03953),
	.w8(32'h3b7e71b2),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b17b79d),
	.w1(32'h3a3402ec),
	.w2(32'hb838ed19),
	.w3(32'h3b5c4f72),
	.w4(32'h3b36782b),
	.w5(32'h3a94a387),
	.w6(32'h3a7ee186),
	.w7(32'h39ba5dae),
	.w8(32'h3a3c78e4),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a756046),
	.w1(32'h3b0d1cd4),
	.w2(32'h3aa95952),
	.w3(32'h3b0cad16),
	.w4(32'h3aa0e553),
	.w5(32'hbb361e62),
	.w6(32'h3aaa1102),
	.w7(32'h3ad21035),
	.w8(32'hbb26cef1),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaba16f9),
	.w1(32'hbafbbf22),
	.w2(32'hbb2c69ef),
	.w3(32'hbb2f7d57),
	.w4(32'hbb17806b),
	.w5(32'hbadce2a5),
	.w6(32'hbb39a2bc),
	.w7(32'hbb416b32),
	.w8(32'hbaf092ce),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba836cf3),
	.w1(32'hb9160e01),
	.w2(32'hb8b4076c),
	.w3(32'hba05af6a),
	.w4(32'hba1e0c88),
	.w5(32'h3980313f),
	.w6(32'hb8f12cfb),
	.w7(32'h388ccf75),
	.w8(32'h3abc2e2e),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7e4315),
	.w1(32'h3b42f8c9),
	.w2(32'h3a036d5c),
	.w3(32'h3af356ad),
	.w4(32'h3b3455ef),
	.w5(32'hbaf02449),
	.w6(32'h3aba12a2),
	.w7(32'h3b0b60f1),
	.w8(32'hb9a865d6),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba841937),
	.w1(32'h3a36c217),
	.w2(32'hba4bb825),
	.w3(32'h388c458c),
	.w4(32'hb8b0e3ba),
	.w5(32'h3bc08c94),
	.w6(32'h3a512c4a),
	.w7(32'hbab434ef),
	.w8(32'h3bdd5bd8),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4eefbe),
	.w1(32'h3b90eeda),
	.w2(32'h3ba526ab),
	.w3(32'h3bd4b8ab),
	.w4(32'h3b92a967),
	.w5(32'h3b012437),
	.w6(32'h3be0e80b),
	.w7(32'h3b568080),
	.w8(32'h3a164914),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d5dba7),
	.w1(32'h3aa256b7),
	.w2(32'h3a6e2077),
	.w3(32'hb6d76233),
	.w4(32'hbb24ce8d),
	.w5(32'h3b030578),
	.w6(32'h3b16e2e4),
	.w7(32'hbab3c433),
	.w8(32'h3b4b8a57),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3accc3d9),
	.w1(32'h3b343901),
	.w2(32'h3b138103),
	.w3(32'h39fc83ce),
	.w4(32'hb9abbe56),
	.w5(32'hbac0704f),
	.w6(32'h3aae6a0b),
	.w7(32'h3a6fd015),
	.w8(32'h394eb198),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afaef05),
	.w1(32'h3afb3748),
	.w2(32'h39f7683b),
	.w3(32'h3a93d54a),
	.w4(32'h3ad232e6),
	.w5(32'h3a6d2c47),
	.w6(32'h3b2e42d5),
	.w7(32'h3ae99051),
	.w8(32'h3a9331f4),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0fc2d1),
	.w1(32'h3a044995),
	.w2(32'hb830e965),
	.w3(32'h3a36a0ff),
	.w4(32'h39974579),
	.w5(32'hba1aaa6d),
	.w6(32'h3b1377cd),
	.w7(32'h3a092e58),
	.w8(32'hbad8379a),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb92ba1a),
	.w1(32'h37dfc1f2),
	.w2(32'h3aa64655),
	.w3(32'hb990f4b1),
	.w4(32'hba71bff7),
	.w5(32'hbb6115e0),
	.w6(32'hba4cf022),
	.w7(32'hbb16a063),
	.w8(32'hbb633f5b),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb221425),
	.w1(32'hb9862aa5),
	.w2(32'hb9277f07),
	.w3(32'hbb143336),
	.w4(32'hbafd53f2),
	.w5(32'hba554e5d),
	.w6(32'hba515e23),
	.w7(32'hba91bdda),
	.w8(32'hb944240b),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacce424),
	.w1(32'hbb946fc6),
	.w2(32'hbb81dec6),
	.w3(32'hbb47db9c),
	.w4(32'hb9dbc033),
	.w5(32'h39efb44f),
	.w6(32'hbb93473c),
	.w7(32'hbb163ef8),
	.w8(32'h3b2bf08d),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5e4d12),
	.w1(32'hb9ce609f),
	.w2(32'hbabfe994),
	.w3(32'h397ca64a),
	.w4(32'h3a5870e4),
	.w5(32'hbb19260e),
	.w6(32'h3af57eac),
	.w7(32'h39679135),
	.w8(32'hbb344f89),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae203ce),
	.w1(32'h3a1e0ce4),
	.w2(32'h3a54a3d2),
	.w3(32'h3aa6ade8),
	.w4(32'h3a92ab81),
	.w5(32'hbb3ed6c4),
	.w6(32'hba8f737c),
	.w7(32'h3a5f0087),
	.w8(32'hba03a911),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3f58c9),
	.w1(32'h3a7f1341),
	.w2(32'h3aec7e1e),
	.w3(32'hbab5f09e),
	.w4(32'h39f3ad51),
	.w5(32'h3b0dc278),
	.w6(32'hba949fcf),
	.w7(32'h3b365431),
	.w8(32'hba17fc2f),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba99e923),
	.w1(32'h3a1adb16),
	.w2(32'h3b2815b3),
	.w3(32'h3b9485b4),
	.w4(32'h3b37647e),
	.w5(32'hbb203fb8),
	.w6(32'h3a2f0bd9),
	.w7(32'h3a9f4028),
	.w8(32'hba6449d6),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a798a48),
	.w1(32'h3b3af4e6),
	.w2(32'h3b2369ea),
	.w3(32'hbac7bbdb),
	.w4(32'hb91060f2),
	.w5(32'h378a6a0d),
	.w6(32'hba97158b),
	.w7(32'h3a82e60b),
	.w8(32'h3a0bac60),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb05b275),
	.w1(32'h3945174f),
	.w2(32'hb942ace8),
	.w3(32'hbb235f7f),
	.w4(32'hbb125b08),
	.w5(32'h3b4ad9e9),
	.w6(32'hb9984517),
	.w7(32'hb9c73892),
	.w8(32'h3b9f86d6),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1137a6),
	.w1(32'h3b902078),
	.w2(32'h3ac10795),
	.w3(32'h3a1bddcd),
	.w4(32'hba08bb19),
	.w5(32'h3ac14ce6),
	.w6(32'h3b685138),
	.w7(32'h391883db),
	.w8(32'h39e6bb38),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b646d18),
	.w1(32'h39c43ba4),
	.w2(32'hba351ff6),
	.w3(32'h3b126b14),
	.w4(32'h3973e9a3),
	.w5(32'hbbbf9963),
	.w6(32'h3af25924),
	.w7(32'h3a5ed6a7),
	.w8(32'hbb7d166c),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule