module layer_8_featuremap_13(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8a0966),
	.w1(32'h3b5e747d),
	.w2(32'h3a2dd86d),
	.w3(32'hbaecacc1),
	.w4(32'h3b60b9c5),
	.w5(32'h3ad072e2),
	.w6(32'h3bf00283),
	.w7(32'hba7b3a2b),
	.w8(32'h3a99e324),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8d03ea),
	.w1(32'hbb36d6fb),
	.w2(32'hbb1ee137),
	.w3(32'hbae87e99),
	.w4(32'hbbebd222),
	.w5(32'hbbe94049),
	.w6(32'h3b04698c),
	.w7(32'hbbc544cc),
	.w8(32'hbb97547f),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9be78c),
	.w1(32'hba760c60),
	.w2(32'hbac2e7c0),
	.w3(32'hbad76e2f),
	.w4(32'hbb8a49ef),
	.w5(32'hbb9dca17),
	.w6(32'hb89c47da),
	.w7(32'hbb4c9fbf),
	.w8(32'hba123f96),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ac5430),
	.w1(32'hbbc2425a),
	.w2(32'hba8b8df2),
	.w3(32'hbbae034b),
	.w4(32'hbbc2b626),
	.w5(32'hbb9307b9),
	.w6(32'h3b06415e),
	.w7(32'hbb791374),
	.w8(32'h3aacd68d),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb04e97f),
	.w1(32'h3b90f3d9),
	.w2(32'h3b0ae19c),
	.w3(32'hbb348de4),
	.w4(32'h3b7ec3f8),
	.w5(32'hbb936cd6),
	.w6(32'h3be5057f),
	.w7(32'h3b72e487),
	.w8(32'h3ba56981),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b90c31b),
	.w1(32'h3b1a5d3d),
	.w2(32'hbbc4f445),
	.w3(32'hbc128b5b),
	.w4(32'h3ac95193),
	.w5(32'h3c8710cb),
	.w6(32'h3b9615d6),
	.w7(32'hbb498fe1),
	.w8(32'hbc8e9824),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb379eee),
	.w1(32'h3a179cfa),
	.w2(32'hb9b710c2),
	.w3(32'hbc154e1c),
	.w4(32'h3ac576ce),
	.w5(32'hba577233),
	.w6(32'h3c5cad5a),
	.w7(32'h3b4cfba9),
	.w8(32'hbaa48c5f),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacd84df),
	.w1(32'h3c1c4f58),
	.w2(32'hbb4c5974),
	.w3(32'h3b2ce7e0),
	.w4(32'hbc0a460c),
	.w5(32'hbb468d02),
	.w6(32'hbbcd59bc),
	.w7(32'hbbae9ac5),
	.w8(32'hbc1acba9),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3270f8),
	.w1(32'h3a9f0ae3),
	.w2(32'hba8cc65b),
	.w3(32'hbbde0279),
	.w4(32'hbb01d8ff),
	.w5(32'hbb3a5375),
	.w6(32'h3a444cbd),
	.w7(32'hbb3995f8),
	.w8(32'hbb3c4b70),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb926e2e),
	.w1(32'hbba8a725),
	.w2(32'h3be7c0be),
	.w3(32'hbbc4dabc),
	.w4(32'hbc1430f4),
	.w5(32'hbc97a39b),
	.w6(32'hbb7025bd),
	.w7(32'h3c944a50),
	.w8(32'h3c520f12),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd5ee4f),
	.w1(32'h3b4c7317),
	.w2(32'hbae43b52),
	.w3(32'h3bad1807),
	.w4(32'h3b5990fc),
	.w5(32'hbbad0810),
	.w6(32'hbc129605),
	.w7(32'hbbb2800d),
	.w8(32'hbba32bd6),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc40fcd9),
	.w1(32'h3abd0f20),
	.w2(32'hba4c3e59),
	.w3(32'hbc276616),
	.w4(32'hbb86d6a9),
	.w5(32'hbb0a9378),
	.w6(32'hbc070fb3),
	.w7(32'h3c1dab30),
	.w8(32'hbc325936),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac0802b),
	.w1(32'h3cabf0a1),
	.w2(32'hbc08a3db),
	.w3(32'hbb366de8),
	.w4(32'hbcf42c6d),
	.w5(32'hbcec4eb6),
	.w6(32'hbb777f5c),
	.w7(32'h3c8c374e),
	.w8(32'h3c7d3bd1),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd3a0692),
	.w1(32'hbbc175c2),
	.w2(32'hbc039600),
	.w3(32'h3d30b092),
	.w4(32'hbb532c64),
	.w5(32'h3b0f38c3),
	.w6(32'hbc972190),
	.w7(32'h38964e2a),
	.w8(32'hbb1ce776),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad8d249),
	.w1(32'h3b6fa97f),
	.w2(32'hba6c33ee),
	.w3(32'hbbd232f9),
	.w4(32'h3b76c043),
	.w5(32'hbb31501e),
	.w6(32'h3b880df9),
	.w7(32'hbafc2f39),
	.w8(32'h3ab34043),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba804edc),
	.w1(32'hbb91a407),
	.w2(32'hbc37ef9c),
	.w3(32'hba9a5c5c),
	.w4(32'h3bc36a6c),
	.w5(32'h3bc4394c),
	.w6(32'hbbbc83fb),
	.w7(32'hbb277a77),
	.w8(32'h3b46e143),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc10e407),
	.w1(32'hbc5c985f),
	.w2(32'hbc59dd42),
	.w3(32'h3b5d1918),
	.w4(32'h3c867a15),
	.w5(32'h3ce00216),
	.w6(32'h3c13f586),
	.w7(32'h3c344c01),
	.w8(32'hbc8094a0),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c541c70),
	.w1(32'h39e33a42),
	.w2(32'hbaeb1407),
	.w3(32'h3be84aaa),
	.w4(32'h3967ebc2),
	.w5(32'h3ad0e2f2),
	.w6(32'hbc853d08),
	.w7(32'hba92eb6c),
	.w8(32'hb9e6721d),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3a4876),
	.w1(32'h3bcbc3ec),
	.w2(32'h3ceb33f8),
	.w3(32'hbac3d435),
	.w4(32'hba360242),
	.w5(32'hbda8bd12),
	.w6(32'hb936265b),
	.w7(32'hbcc6aa41),
	.w8(32'h3d3e0d70),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbce8d545),
	.w1(32'h3b9c0618),
	.w2(32'h3ae526cc),
	.w3(32'hbbe37331),
	.w4(32'h3ba299cc),
	.w5(32'hbb804ca0),
	.w6(32'h3c3c5e58),
	.w7(32'h3b3b0ed1),
	.w8(32'h3a2e93ec),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb3f26e),
	.w1(32'hbb9c0264),
	.w2(32'hbbddaaaa),
	.w3(32'hbaad9376),
	.w4(32'hbb0d8386),
	.w5(32'h3b25794c),
	.w6(32'hbbaf51aa),
	.w7(32'hbb580b2c),
	.w8(32'hbb167d91),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5464cf),
	.w1(32'hbc33fa71),
	.w2(32'h3c0293f6),
	.w3(32'hba84395d),
	.w4(32'h3cd989fc),
	.w5(32'hbb924962),
	.w6(32'h3b47c2ba),
	.w7(32'hbd0426d1),
	.w8(32'hba5530f6),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c18d845),
	.w1(32'h3cbf8036),
	.w2(32'hbc801082),
	.w3(32'hbb860536),
	.w4(32'hbd2fefac),
	.w5(32'h3cfd87d7),
	.w6(32'hbc81ecc1),
	.w7(32'h3cff36b9),
	.w8(32'hbb8a3297),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc177e29),
	.w1(32'h3b07b9bd),
	.w2(32'hbaa17850),
	.w3(32'h3cdff710),
	.w4(32'h3b04478c),
	.w5(32'hbaa188a8),
	.w6(32'hbd26c66b),
	.w7(32'h3a200b5d),
	.w8(32'hbb0c627c),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb29f3f1),
	.w1(32'hbc0323ef),
	.w2(32'hb998b495),
	.w3(32'h3b44d2ab),
	.w4(32'hbbd6ac36),
	.w5(32'hbd13d321),
	.w6(32'hbb522b67),
	.w7(32'hbcc050f3),
	.w8(32'hbaf7a31b),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca893bd),
	.w1(32'h3ba8ba64),
	.w2(32'h3ad8956f),
	.w3(32'hbabf54ab),
	.w4(32'hbb4c08e7),
	.w5(32'h3b74756a),
	.w6(32'hbcf8d9dc),
	.w7(32'h3bf34789),
	.w8(32'h3b04f2e7),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc027627),
	.w1(32'h3aab3c3a),
	.w2(32'hbbb17436),
	.w3(32'h3b4d8788),
	.w4(32'h3b50e039),
	.w5(32'h3b5fc0fd),
	.w6(32'hbc330c0b),
	.w7(32'hbb68c096),
	.w8(32'hbb05f3f8),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4c452f),
	.w1(32'hbc525dc1),
	.w2(32'hbc66c048),
	.w3(32'h3adc6a08),
	.w4(32'hbc5b2a5a),
	.w5(32'hbc8af6c2),
	.w6(32'h3822859a),
	.w7(32'hbbbd8bc7),
	.w8(32'hbc1aabb0),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7bd74c),
	.w1(32'h3b267357),
	.w2(32'hbb45e123),
	.w3(32'h3b73d308),
	.w4(32'h3b81bfd2),
	.w5(32'h3b320550),
	.w6(32'hbc28337f),
	.w7(32'hbbaa5cd8),
	.w8(32'h39f85a95),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7af264),
	.w1(32'h3aefeb30),
	.w2(32'hbb2c31f8),
	.w3(32'hbbdead8b),
	.w4(32'h3b57ea48),
	.w5(32'h3b5c8085),
	.w6(32'h3b04b7fe),
	.w7(32'hb95a09cb),
	.w8(32'hbb6812c6),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb755fb0),
	.w1(32'hbb883d47),
	.w2(32'hbc812d1f),
	.w3(32'hba5712f3),
	.w4(32'hbb882db0),
	.w5(32'hbcb7ae75),
	.w6(32'hbb1585ee),
	.w7(32'hbb87ae6d),
	.w8(32'hbc862581),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3cfa8d),
	.w1(32'h3b8543be),
	.w2(32'h3af81c56),
	.w3(32'hbc78b909),
	.w4(32'hb93c589f),
	.w5(32'h3aff1eaf),
	.w6(32'h3b23d108),
	.w7(32'hbb2d150e),
	.w8(32'hbbca6e56),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b56b026),
	.w1(32'h3a86c94f),
	.w2(32'h3ae39d6c),
	.w3(32'h3a7d69d0),
	.w4(32'h3b322e66),
	.w5(32'hb946c720),
	.w6(32'hb9d4dd5e),
	.w7(32'h3b63a4b2),
	.w8(32'h3b076b0a),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1dd212),
	.w1(32'h3a93e493),
	.w2(32'h3bbd3577),
	.w3(32'h39df8556),
	.w4(32'h3c6bb2b4),
	.w5(32'hbc91f88a),
	.w6(32'h3ad081f1),
	.w7(32'hbc0855f3),
	.w8(32'hbbfd2994),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3fe09c),
	.w1(32'h3b379d53),
	.w2(32'h3ab9206f),
	.w3(32'hbba6dae1),
	.w4(32'h3a2dfa5e),
	.w5(32'h3b03f136),
	.w6(32'h3ab78f5e),
	.w7(32'h3a80357c),
	.w8(32'h3a875136),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba59256),
	.w1(32'hbb3794ed),
	.w2(32'hbb9213ec),
	.w3(32'h391a60c0),
	.w4(32'hbc1fd741),
	.w5(32'hbb3d2579),
	.w6(32'h3b8437f8),
	.w7(32'hbc2fb662),
	.w8(32'hbb7fcd50),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4e841e),
	.w1(32'hbb25338e),
	.w2(32'hbc8ecb1d),
	.w3(32'hbb1911a2),
	.w4(32'hbc201fe1),
	.w5(32'h3aee91c9),
	.w6(32'h3b990f13),
	.w7(32'h3c583336),
	.w8(32'hbc08dd7e),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcaa06ac),
	.w1(32'hbc2814b4),
	.w2(32'hbc729c84),
	.w3(32'h3c86de86),
	.w4(32'h3b95a53f),
	.w5(32'h3c1cbb03),
	.w6(32'hbc0e0e8f),
	.w7(32'h3bc44678),
	.w8(32'hbbeb0439),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4759d3),
	.w1(32'hbc60efc1),
	.w2(32'h3ba5a96d),
	.w3(32'h3a66dd99),
	.w4(32'hbd1398e8),
	.w5(32'hbcffada9),
	.w6(32'hbc1cd756),
	.w7(32'hbc54e600),
	.w8(32'hbbab7941),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0d544e),
	.w1(32'hbba872df),
	.w2(32'hbbe9d5b0),
	.w3(32'hbd377a13),
	.w4(32'hbb6571ae),
	.w5(32'hbb8bfee9),
	.w6(32'hbc91decb),
	.w7(32'h39d1c612),
	.w8(32'hbbff8f57),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39858bac),
	.w1(32'hbbb38a2f),
	.w2(32'h3ae78a78),
	.w3(32'hbb94b260),
	.w4(32'h3beeb8cc),
	.w5(32'h3c746779),
	.w6(32'hb96d0989),
	.w7(32'h3c120556),
	.w8(32'h3c54960f),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdfd53f),
	.w1(32'hbb1cc044),
	.w2(32'hbb28836f),
	.w3(32'h3c79c76e),
	.w4(32'h3af16e7a),
	.w5(32'h3aec21c6),
	.w6(32'h3b5918ae),
	.w7(32'h3b49a660),
	.w8(32'h3b185203),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab4b079),
	.w1(32'h3b0b053b),
	.w2(32'h3b4f92fe),
	.w3(32'hbb628317),
	.w4(32'h3b7a5426),
	.w5(32'h3b5fab2a),
	.w6(32'h3ba92346),
	.w7(32'h3b30867b),
	.w8(32'h3b3efba0),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6d0aff),
	.w1(32'hbb6a3cc1),
	.w2(32'hbbd95526),
	.w3(32'h3afb1c30),
	.w4(32'h3b4fcb97),
	.w5(32'hbc224dca),
	.w6(32'h3a512431),
	.w7(32'h3a047057),
	.w8(32'hbc3896b3),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0f5d60),
	.w1(32'hbcdeea88),
	.w2(32'hbb388fbd),
	.w3(32'hbbbc01b2),
	.w4(32'h3cc6a240),
	.w5(32'h3cf7c519),
	.w6(32'hbcb0f599),
	.w7(32'hbbb52655),
	.w8(32'hbca73456),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d0c5b90),
	.w1(32'hbba0da4d),
	.w2(32'h3ab11e87),
	.w3(32'hbce27f57),
	.w4(32'h3c4d43d1),
	.w5(32'hbb969b7f),
	.w6(32'h3cdbfdc0),
	.w7(32'hbc60e66b),
	.w8(32'hbc935e3f),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc015ac),
	.w1(32'h3c594410),
	.w2(32'hbc9f5285),
	.w3(32'hbc6f678a),
	.w4(32'hbb986284),
	.w5(32'h3ba3338e),
	.w6(32'hbc8bfa77),
	.w7(32'hbc8a761f),
	.w8(32'hbcb60deb),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8aa2cc),
	.w1(32'hbb2bb0ec),
	.w2(32'hbbddd6dc),
	.w3(32'hbcc1f19b),
	.w4(32'hbccaac7d),
	.w5(32'hbc80fb26),
	.w6(32'h3c14392e),
	.w7(32'hbb7282ae),
	.w8(32'hbb9d81e9),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc093ee1),
	.w1(32'h3c00ee88),
	.w2(32'h3b6db801),
	.w3(32'hbcc3acee),
	.w4(32'h39f6880e),
	.w5(32'hbae1a352),
	.w6(32'hba7f88e8),
	.w7(32'h37207945),
	.w8(32'h3a25d75b),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a921e4e),
	.w1(32'h3c1e35ea),
	.w2(32'h3b1c4316),
	.w3(32'h3a832e8d),
	.w4(32'hbb86a28e),
	.w5(32'hbb6261ee),
	.w6(32'hbbc2c10a),
	.w7(32'hba0fee9c),
	.w8(32'h3c23add8),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbce5bdd),
	.w1(32'hba69f9b7),
	.w2(32'hb854fedb),
	.w3(32'h3b454c13),
	.w4(32'h3a2c3e57),
	.w5(32'hbb9734ce),
	.w6(32'h3b6511f1),
	.w7(32'hbae34512),
	.w8(32'h3ad8949d),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b842017),
	.w1(32'h39b71fa3),
	.w2(32'h3a9bc1c0),
	.w3(32'hbb21e897),
	.w4(32'h3a913e81),
	.w5(32'hbaff42b0),
	.w6(32'hbbf65cc1),
	.w7(32'h3a74762f),
	.w8(32'h3acef9fb),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b211ee9),
	.w1(32'hbc30e17d),
	.w2(32'hbbc48d63),
	.w3(32'h396ac360),
	.w4(32'h3ce589f6),
	.w5(32'h3d2ffeb3),
	.w6(32'h3b5950fc),
	.w7(32'h3c1bd987),
	.w8(32'h3c04b94f),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cf105e3),
	.w1(32'h3ad90141),
	.w2(32'h3d0ea40c),
	.w3(32'hbc0bb8e7),
	.w4(32'h3d19dbdc),
	.w5(32'hbd4ff150),
	.w6(32'h3d08ab01),
	.w7(32'hbd31ce6c),
	.w8(32'h3d0ace3a),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6b85f3),
	.w1(32'hbb996e6d),
	.w2(32'h3c98c515),
	.w3(32'hbd49d8e8),
	.w4(32'h3ccee527),
	.w5(32'h3c357de3),
	.w6(32'h3d35d602),
	.w7(32'hbcc36fa1),
	.w8(32'hbc294d89),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d365cc3),
	.w1(32'h3a9836e2),
	.w2(32'hbaac98d4),
	.w3(32'hbd0c3ecb),
	.w4(32'h3aa493aa),
	.w5(32'h39e0a47c),
	.w6(32'hba378a5a),
	.w7(32'h3a07f820),
	.w8(32'hba1f2e87),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d6ba2b),
	.w1(32'hba4085dc),
	.w2(32'h3b3be071),
	.w3(32'hba09e1dd),
	.w4(32'h3b5321b0),
	.w5(32'h3ab16c2f),
	.w6(32'h3a90b749),
	.w7(32'hbaafb973),
	.w8(32'h3ba9e045),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbdaabd),
	.w1(32'hbbdbe71f),
	.w2(32'h3a212d6e),
	.w3(32'hb883e612),
	.w4(32'h3a7eaeea),
	.w5(32'hbbac4a2b),
	.w6(32'hbc189885),
	.w7(32'hbb3c1b14),
	.w8(32'hbbf3080b),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe81e9c),
	.w1(32'hbb05c30d),
	.w2(32'hbab4aab9),
	.w3(32'hbb93dac6),
	.w4(32'hbaf5646a),
	.w5(32'h3aa1435b),
	.w6(32'hbc8984c6),
	.w7(32'hba08d104),
	.w8(32'h399d3640),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3075ce),
	.w1(32'hbb73a128),
	.w2(32'h3d0d542f),
	.w3(32'h396aaf55),
	.w4(32'h3c194910),
	.w5(32'h3889434b),
	.w6(32'hbb97ff9d),
	.w7(32'h3cb12170),
	.w8(32'h3d02924f),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7322b0),
	.w1(32'hba444ccd),
	.w2(32'hbbb41171),
	.w3(32'h3d28179e),
	.w4(32'h3b785944),
	.w5(32'hba05705d),
	.w6(32'hbcd12143),
	.w7(32'h3ac180d4),
	.w8(32'h3ad95cce),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc8feff),
	.w1(32'h3bd518b6),
	.w2(32'hbc9ed3dd),
	.w3(32'hbb1015d3),
	.w4(32'hbbead303),
	.w5(32'hbaf26589),
	.w6(32'h3c6d372f),
	.w7(32'hbb8dccd6),
	.w8(32'hbc82f2d1),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0bee67),
	.w1(32'h3b374cf2),
	.w2(32'hbb2ed719),
	.w3(32'h3b77ee49),
	.w4(32'hba020a84),
	.w5(32'hbb64d0b6),
	.w6(32'h3c1e2836),
	.w7(32'hba365bbe),
	.w8(32'hbb05f0ba),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf16213),
	.w1(32'hbaefb20d),
	.w2(32'h3ceec872),
	.w3(32'hbbd308b8),
	.w4(32'h3d16a088),
	.w5(32'hbd49546c),
	.w6(32'hbae63767),
	.w7(32'hbd52dcf5),
	.w8(32'h3cbe1eb2),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c216fbf),
	.w1(32'h3b3071a8),
	.w2(32'hbb96d392),
	.w3(32'hbd3ccbeb),
	.w4(32'h3b0a9608),
	.w5(32'h3b243527),
	.w6(32'h3d328551),
	.w7(32'h3adb5407),
	.w8(32'hb8cd8634),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb65d1b5),
	.w1(32'hba876f39),
	.w2(32'hb866ca90),
	.w3(32'h3aead0f2),
	.w4(32'h3a8020c5),
	.w5(32'h3b901f31),
	.w6(32'h3987f024),
	.w7(32'h3ae3f5cd),
	.w8(32'h3ba1eef7),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc604aa),
	.w1(32'hbb982f74),
	.w2(32'hbbfb8f00),
	.w3(32'h3bf4da5f),
	.w4(32'hbb7fdf57),
	.w5(32'h3a47c3c4),
	.w6(32'h3bd444ad),
	.w7(32'hbbc7f218),
	.w8(32'hbbcda9d8),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb178142),
	.w1(32'hbb7a483c),
	.w2(32'hbbe6c09d),
	.w3(32'hbc08e9ee),
	.w4(32'h3936b544),
	.w5(32'h3c0f208f),
	.w6(32'hbabdb2ea),
	.w7(32'h38e143a2),
	.w8(32'hb9c06cef),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a1cf3),
	.w1(32'h3a64818c),
	.w2(32'hbb6593d6),
	.w3(32'hbb7edb12),
	.w4(32'h3abc1ff5),
	.w5(32'h3bb5a4e4),
	.w6(32'h3b63a554),
	.w7(32'h3b136038),
	.w8(32'hba9bdb8a),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc09daa5),
	.w1(32'hbf3c34a8),
	.w2(32'hbea6ffff),
	.w3(32'h3b638312),
	.w4(32'hbf3011fc),
	.w5(32'hbef095bf),
	.w6(32'hbb36015f),
	.w7(32'hbfc014a7),
	.w8(32'hbf5e8740),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbeb5138a),
	.w1(32'hbf921f83),
	.w2(32'hbe7de382),
	.w3(32'h3f8c3bc3),
	.w4(32'hc01961c6),
	.w5(32'hbf38d55e),
	.w6(32'hbecc3d8b),
	.w7(32'hbf2582e3),
	.w8(32'hbf65bf23),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbf61579d),
	.w1(32'hbf237276),
	.w2(32'hbe32a222),
	.w3(32'hbf60c94e),
	.w4(32'hbf3fc0c2),
	.w5(32'hbf13bd82),
	.w6(32'h3fbfede4),
	.w7(32'hbee869b1),
	.w8(32'hbf3408bc),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbf530a12),
	.w1(32'hbe9864e8),
	.w2(32'hbebf8e62),
	.w3(32'hbf370258),
	.w4(32'h3fa9f00c),
	.w5(32'hbf814d32),
	.w6(32'hbf027253),
	.w7(32'hbf4b89b3),
	.w8(32'hbf13f644),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbf495852),
	.w1(32'h3fe2711c),
	.w2(32'hbf56eb3c),
	.w3(32'hbf87fe65),
	.w4(32'h3ef79733),
	.w5(32'hbf217482),
	.w6(32'hbf380c13),
	.w7(32'hbf2eec5d),
	.w8(32'hbf1a3a73),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbf242efd),
	.w1(32'h3fbae543),
	.w2(32'h3fae3ef8),
	.w3(32'hbef072f5),
	.w4(32'hbf17fac7),
	.w5(32'h3f948d08),
	.w6(32'hbe9ff6ee),
	.w7(32'hbf03d817),
	.w8(32'hbebd70dc),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbf26afcc),
	.w1(32'hbfac9ee6),
	.w2(32'h3fc54012),
	.w3(32'hbf55bf09),
	.w4(32'hbf2106fc),
	.w5(32'hbf35f3a7),
	.w6(32'hbf3021c6),
	.w7(32'hbf3d6806),
	.w8(32'hbee63642),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbf9ae113),
	.w1(32'h3ef391da),
	.w2(32'h3f4b2f2b),
	.w3(32'h3f3a4017),
	.w4(32'h3ee83a30),
	.w5(32'h3ebef258),
	.w6(32'hbf0e2db1),
	.w7(32'h3f3a1e47),
	.w8(32'h3edbe91f),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f5180b6),
	.w1(32'h3ed70447),
	.w2(32'h3f4a2d2f),
	.w3(32'h3ed49444),
	.w4(32'h3f16963b),
	.w5(32'h3f0d8c44),
	.w6(32'h3e9ab073),
	.w7(32'h3fa1f7a0),
	.w8(32'h3f4b9b16),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f20a428),
	.w1(32'h3da9811b),
	.w2(32'h3ef06c08),
	.w3(32'h3f08879a),
	.w4(32'h3f1d37ba),
	.w5(32'h3eb4c2c9),
	.w6(32'h3f337650),
	.w7(32'h3f463944),
	.w8(32'h3f3f5508),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3edb15b6),
	.w1(32'h3ef328e5),
	.w2(32'h3ef1c9e1),
	.w3(32'h3ee42898),
	.w4(32'h3ea57487),
	.w5(32'h3ec17c33),
	.w6(32'h3ecca170),
	.w7(32'h3ed99201),
	.w8(32'h3f1d4870),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f291e8c),
	.w1(32'h3ef0713b),
	.w2(32'h3eb4c446),
	.w3(32'h3f152dae),
	.w4(32'h3ef2938a),
	.w5(32'h3f65d474),
	.w6(32'h3f12f945),
	.w7(32'h3e8fb315),
	.w8(32'h3ed38162),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f16fa2d),
	.w1(32'h3ec4131a),
	.w2(32'h3f21b7f8),
	.w3(32'h3f4c715f),
	.w4(32'h3ecc9cbd),
	.w5(32'h3ebf8458),
	.w6(32'h3f0cbdf0),
	.w7(32'h3ee91143),
	.w8(32'h3ea3db80),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f0af726),
	.w1(32'h3f2fca59),
	.w2(32'h3f294de0),
	.w3(32'h3f3b0912),
	.w4(32'h3fa0b576),
	.w5(32'h3ed49eb1),
	.w6(32'h3edbdab2),
	.w7(32'h3f4abd4f),
	.w8(32'h3f00925a),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f26cf64),
	.w1(32'h3f2864f0),
	.w2(32'hbde83fd3),
	.w3(32'h3f22057d),
	.w4(32'h3e1fca21),
	.w5(32'h3da85436),
	.w6(32'h3f03b04e),
	.w7(32'h3dd53ec3),
	.w8(32'h3ce91754),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9328cd),
	.w1(32'h3b75a8bb),
	.w2(32'h3d7d5052),
	.w3(32'hbdeaf44e),
	.w4(32'h3d027b2e),
	.w5(32'hbe5d53ef),
	.w6(32'h3c95a633),
	.w7(32'h3bd333bb),
	.w8(32'hbce92505),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbe8e5ae6),
	.w1(32'hbdecbf77),
	.w2(32'hbe2089b2),
	.w3(32'h3c20e606),
	.w4(32'h3ddd0100),
	.w5(32'h3d638d6d),
	.w6(32'h3c12c7b0),
	.w7(32'h3d97e094),
	.w8(32'hbc52e248),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbdc61b1b),
	.w1(32'h3c476303),
	.w2(32'h3db4f22f),
	.w3(32'h3dd77b09),
	.w4(32'hbd177c93),
	.w5(32'h3dacad45),
	.w6(32'h3d3b6cf1),
	.w7(32'h3c8b7e2b),
	.w8(32'h3cf5577c),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3da3b883),
	.w1(32'h3d863c7b),
	.w2(32'h3d41c72b),
	.w3(32'hbe293d4a),
	.w4(32'h3d8ada86),
	.w5(32'h3d97bcb8),
	.w6(32'h3d57af9b),
	.w7(32'h3dde1c1f),
	.w8(32'hbe413410),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d8116cd),
	.w1(32'hbcc4ee3a),
	.w2(32'h3e01a621),
	.w3(32'hbc4ed068),
	.w4(32'h3c09df1a),
	.w5(32'h3e20fa7a),
	.w6(32'hbe1840ac),
	.w7(32'h3be39d4a),
	.w8(32'h3bcff96c),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baef961),
	.w1(32'h3c7657aa),
	.w2(32'h3e0bf085),
	.w3(32'hbcb1c150),
	.w4(32'hbdd303a1),
	.w5(32'hbd7a2d06),
	.w6(32'hbdeb76a4),
	.w7(32'h3e32b01f),
	.w8(32'h3dc1d05e),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3dcaf09d),
	.w1(32'h3de27c9b),
	.w2(32'h3b7743c3),
	.w3(32'h3d16dac2),
	.w4(32'h3d9bf194),
	.w5(32'h3d11f5b6),
	.w6(32'h3bb86f69),
	.w7(32'hb9203334),
	.w8(32'h3cb0c8cc),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cae5173),
	.w1(32'h3c24589e),
	.w2(32'h3bfeae8e),
	.w3(32'h3becdcef),
	.w4(32'h3e5f84ba),
	.w5(32'h3d338cb6),
	.w6(32'h3cdb51e7),
	.w7(32'h3cfdf222),
	.w8(32'h3d1e0994),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3dcb7693),
	.w1(32'h3c0bd554),
	.w2(32'h3c8ec69a),
	.w3(32'h3d01143e),
	.w4(32'h3cd61495),
	.w5(32'h3cca30e5),
	.w6(32'h3c387c58),
	.w7(32'h3b9ba41b),
	.w8(32'h3c64e6ab),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d024893),
	.w1(32'h3baf7c85),
	.w2(32'h3c817663),
	.w3(32'h3d2456dd),
	.w4(32'h3b65410f),
	.w5(32'h3ee02d54),
	.w6(32'h3b156e8a),
	.w7(32'h3bfab050),
	.w8(32'h3b4b9799),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca0c074),
	.w1(32'h3c78e387),
	.w2(32'h3f0a1b6a),
	.w3(32'h3bb8f824),
	.w4(32'h3c2b5bc7),
	.w5(32'h3e3f8a4b),
	.w6(32'h3cf2a84b),
	.w7(32'h3c0db612),
	.w8(32'h3b3cc760),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d0a3a02),
	.w1(32'h3d1e90aa),
	.w2(32'h3ec3b473),
	.w3(32'h3b690925),
	.w4(32'h3d1976e2),
	.w5(32'h3b98e7b8),
	.w6(32'h3cb0d573),
	.w7(32'h3ce4c3ff),
	.w8(32'h3d003553),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3eaafe22),
	.w1(32'h3cfecaec),
	.w2(32'h3dd4fa17),
	.w3(32'h3e7a168e),
	.w4(32'h3b89f879),
	.w5(32'h3d0c47b0),
	.w6(32'h3d7c81db),
	.w7(32'h3cdf2a76),
	.w8(32'h3c81ad0e),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ed4d817),
	.w1(32'h3bd10b94),
	.w2(32'h3d71ab84),
	.w3(32'h3c2cb1c2),
	.w4(32'h3f09ca1d),
	.w5(32'hba58ca04),
	.w6(32'h3d3ca487),
	.w7(32'h3d8f9ebf),
	.w8(32'h3ad2df6e),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb441974),
	.w1(32'h3c873acd),
	.w2(32'h3b6a59af),
	.w3(32'h3bc3b1ed),
	.w4(32'h3bab41d9),
	.w5(32'hbb2eefdb),
	.w6(32'hba199aef),
	.w7(32'hbbb4f558),
	.w8(32'h3c295b15),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afd806b),
	.w1(32'h3c0fe413),
	.w2(32'hb94c8a5d),
	.w3(32'h3b90856d),
	.w4(32'hbaec2325),
	.w5(32'h379fc735),
	.w6(32'h399ca9eb),
	.w7(32'h3c2febc8),
	.w8(32'hbb6e060b),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0a2d45),
	.w1(32'hbb849d42),
	.w2(32'h3b40aca4),
	.w3(32'h3adfcd70),
	.w4(32'hbbb9d30d),
	.w5(32'h392c94f6),
	.w6(32'hbb75c37d),
	.w7(32'hbaf0936b),
	.w8(32'h3a53c503),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd17d9f),
	.w1(32'h3aa3cdf6),
	.w2(32'h3aab4213),
	.w3(32'hbaf2ec96),
	.w4(32'h3b98fe0f),
	.w5(32'h3adb91d0),
	.w6(32'h3aa25c4e),
	.w7(32'h3bd7d01e),
	.w8(32'hbb3905c0),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a150ccf),
	.w1(32'hb959aa0a),
	.w2(32'h3ae2b7e2),
	.w3(32'h3bbf45c7),
	.w4(32'hba36e5d9),
	.w5(32'hbb8a23e0),
	.w6(32'hbbb3ea98),
	.w7(32'hbb0f3cd2),
	.w8(32'h3c2e95fd),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb023eb2),
	.w1(32'hbba77bd6),
	.w2(32'hb888b9d0),
	.w3(32'h3c3bdeff),
	.w4(32'hbb856e26),
	.w5(32'h3980a0d8),
	.w6(32'hbb631d2f),
	.w7(32'hba9b0189),
	.w8(32'h3a179d43),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37b8d178),
	.w1(32'h3a1cfd39),
	.w2(32'h3bf25ddf),
	.w3(32'hbae8a656),
	.w4(32'h3b572541),
	.w5(32'h3b9847a9),
	.w6(32'h38a984e2),
	.w7(32'hbb8d7fc5),
	.w8(32'hbb915655),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0e6035),
	.w1(32'h3bd0c8b2),
	.w2(32'hba07944e),
	.w3(32'h3aa55a3b),
	.w4(32'hbbd0fe81),
	.w5(32'h3b0f0f05),
	.w6(32'hba3c6933),
	.w7(32'hbb03e3f3),
	.w8(32'h3b151355),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb462061),
	.w1(32'hbb93310a),
	.w2(32'h3c8c9bc9),
	.w3(32'h3ba1b026),
	.w4(32'h3ac8565e),
	.w5(32'hbba04fcd),
	.w6(32'h3ace2a57),
	.w7(32'h3bb107d5),
	.w8(32'hbbdb0792),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h388c6bd9),
	.w1(32'h3bd64e97),
	.w2(32'hba232482),
	.w3(32'h3af60ec1),
	.w4(32'h3b90cefc),
	.w5(32'h38f3508f),
	.w6(32'hba8893bf),
	.w7(32'h394f9182),
	.w8(32'hbba70ee7),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0f27ae),
	.w1(32'hba9e8ba5),
	.w2(32'hbb3e3501),
	.w3(32'h3c04539d),
	.w4(32'hbaaf2d64),
	.w5(32'hbc08a195),
	.w6(32'hbb482c80),
	.w7(32'h39dd49aa),
	.w8(32'hbbed7d09),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa4aff7),
	.w1(32'hbaea960c),
	.w2(32'h3b16c34f),
	.w3(32'h3c02adec),
	.w4(32'h3beae575),
	.w5(32'h3c5b4196),
	.w6(32'h3b7a2949),
	.w7(32'hbb72e44b),
	.w8(32'h3c3783e2),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba39fe67),
	.w1(32'h3b6d0a72),
	.w2(32'h3ad61e98),
	.w3(32'hbbba8eba),
	.w4(32'h3bd95510),
	.w5(32'hbb3ef97b),
	.w6(32'hbb488834),
	.w7(32'hbb3cddc1),
	.w8(32'hbb8effa0),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb6b508),
	.w1(32'hba352e67),
	.w2(32'h3b58f642),
	.w3(32'hbae8d266),
	.w4(32'h3aa0c074),
	.w5(32'h3c0f8423),
	.w6(32'hb9cd92f6),
	.w7(32'hbb2ad638),
	.w8(32'hbbd58d69),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbab5b23),
	.w1(32'h3b63c4bf),
	.w2(32'hbbf98510),
	.w3(32'h3ca45358),
	.w4(32'hbc2d7d7d),
	.w5(32'h3d4ae3d7),
	.w6(32'hbbc55f10),
	.w7(32'h3c0a160a),
	.w8(32'hbbb71e2f),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc283afe),
	.w1(32'h3c324947),
	.w2(32'hbc946991),
	.w3(32'hbb15ee9d),
	.w4(32'h3cf06f6f),
	.w5(32'hbaa17a45),
	.w6(32'hbd20b3c9),
	.w7(32'h3bf60197),
	.w8(32'h3c0055d2),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeabcfa),
	.w1(32'h39e34c40),
	.w2(32'hbcaabdc0),
	.w3(32'h3ca2b26c),
	.w4(32'hbc85b126),
	.w5(32'hbc891f78),
	.w6(32'h3cd59065),
	.w7(32'hbc4e18ad),
	.w8(32'h3b52f819),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcccbd20),
	.w1(32'h3cdd73c4),
	.w2(32'h3bdf4f7c),
	.w3(32'hbbb73517),
	.w4(32'hbc508e93),
	.w5(32'hbce7c188),
	.w6(32'h3cadf081),
	.w7(32'hbbab5d94),
	.w8(32'h3bd2abd2),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd4d1db),
	.w1(32'hba6e3101),
	.w2(32'h3bc50e09),
	.w3(32'hbb3ab8f5),
	.w4(32'hba9b6bf4),
	.w5(32'hbd23961a),
	.w6(32'h3a88eb89),
	.w7(32'hbc2f5565),
	.w8(32'h3c8a818c),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cd5db2b),
	.w1(32'hbca3d83b),
	.w2(32'h3da3fd3e),
	.w3(32'hbd4d1da8),
	.w4(32'hbc04234d),
	.w5(32'h3b8654fe),
	.w6(32'hbb7d91e0),
	.w7(32'hbc0d7e5f),
	.w8(32'h3cbca083),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb98f912),
	.w1(32'h3bcbc7e5),
	.w2(32'h3ba3cbf3),
	.w3(32'h3ac23ef0),
	.w4(32'h3c73bb62),
	.w5(32'hbc10cebc),
	.w6(32'hbca4c007),
	.w7(32'h39e7bc34),
	.w8(32'hbb80385a),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3f3ff5),
	.w1(32'h3c483ce7),
	.w2(32'hbc7180a7),
	.w3(32'h3c11e7f7),
	.w4(32'hbc91842f),
	.w5(32'hbc5968e3),
	.w6(32'h3bd0e0d0),
	.w7(32'hbc8d0882),
	.w8(32'hbc8f19e3),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc52e62),
	.w1(32'hbd02a062),
	.w2(32'h3ad9debe),
	.w3(32'hbc109363),
	.w4(32'hba8468ba),
	.w5(32'h3c92be35),
	.w6(32'hbaed8cca),
	.w7(32'hbc5030e5),
	.w8(32'h3ac5fd1f),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc877016),
	.w1(32'h3c79adf4),
	.w2(32'hbc01ff47),
	.w3(32'hbbc502e8),
	.w4(32'hbbec4ecd),
	.w5(32'hba0d2c95),
	.w6(32'hbc080fe7),
	.w7(32'hbc52b1d6),
	.w8(32'h3c0723cf),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3837b3a1),
	.w1(32'hbc134e29),
	.w2(32'h3d4e0d12),
	.w3(32'hbcfa13d1),
	.w4(32'h3b919087),
	.w5(32'h3a811b5e),
	.w6(32'h3beb2e53),
	.w7(32'hbb4934d8),
	.w8(32'h3c3a2f7e),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9e9686),
	.w1(32'hbc8e3fa1),
	.w2(32'hbc030fb9),
	.w3(32'h3c2e24a8),
	.w4(32'hbc2282e5),
	.w5(32'hbb75ccb6),
	.w6(32'hbb8260ec),
	.w7(32'hbbddd150),
	.w8(32'h3a5cf48b),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a311ee8),
	.w1(32'hbc20614d),
	.w2(32'h3c6e6721),
	.w3(32'h3aac3fa2),
	.w4(32'hbc05d09e),
	.w5(32'hbb0fab1b),
	.w6(32'hbb83aeba),
	.w7(32'h3bab75cb),
	.w8(32'h3b0c4295),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h390d1a0f),
	.w1(32'hbcae6247),
	.w2(32'h3b5ec0ab),
	.w3(32'h3c159540),
	.w4(32'hbac75e5c),
	.w5(32'h3b9e6460),
	.w6(32'h3c66e490),
	.w7(32'hbb5e11ee),
	.w8(32'h3c167af4),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb816cb4),
	.w1(32'h3c029af2),
	.w2(32'hbb835968),
	.w3(32'hbc60c490),
	.w4(32'h3a8eb756),
	.w5(32'h39fdd764),
	.w6(32'h3a9c3f19),
	.w7(32'h3bd03678),
	.w8(32'h3bea1eb1),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb58efbb),
	.w1(32'h3cc12b2c),
	.w2(32'hbb6c38c7),
	.w3(32'hb8f86ef3),
	.w4(32'h3c109182),
	.w5(32'h3bfcde9f),
	.w6(32'hb97f332e),
	.w7(32'h3a9f44d8),
	.w8(32'hbb027012),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule