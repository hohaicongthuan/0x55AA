module layer_10_featuremap_378(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9351139),
	.w1(32'h3b4b8b1f),
	.w2(32'hbc2cd5ff),
	.w3(32'h3c089fa8),
	.w4(32'h3babe0de),
	.w5(32'h3c2ac731),
	.w6(32'h3c2e3b5f),
	.w7(32'hbc938dd5),
	.w8(32'hba20626b),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc901e3e),
	.w1(32'hbba8b03f),
	.w2(32'hbc2a23c5),
	.w3(32'hbb27057b),
	.w4(32'h3bad7052),
	.w5(32'hbb948c58),
	.w6(32'h3b7b32bd),
	.w7(32'hbc4d00b8),
	.w8(32'h3bb753ba),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2d85c4),
	.w1(32'hbbc09f80),
	.w2(32'h3b908265),
	.w3(32'hbc9dd6f5),
	.w4(32'hbcc595cb),
	.w5(32'hb991e5d7),
	.w6(32'h3bec0414),
	.w7(32'hbbc4424a),
	.w8(32'h3a465c3e),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b801ea9),
	.w1(32'hbbea4cc6),
	.w2(32'h3bb37ef7),
	.w3(32'hbc4f4539),
	.w4(32'hbc0d2a0d),
	.w5(32'hbbc8789b),
	.w6(32'h3bd992e3),
	.w7(32'h3a85b276),
	.w8(32'hbc14c681),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0fba46),
	.w1(32'hba9e52d4),
	.w2(32'hbb5dc903),
	.w3(32'hbb5622d8),
	.w4(32'h3b4b55be),
	.w5(32'hba3140b9),
	.w6(32'h3b2ee01c),
	.w7(32'h3a35f30b),
	.w8(32'hba348cbd),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3a7595),
	.w1(32'hbc24033a),
	.w2(32'h3a929158),
	.w3(32'hbc193b86),
	.w4(32'hbaeb43c7),
	.w5(32'hbab37f7b),
	.w6(32'h3b9a533f),
	.w7(32'h3c52748f),
	.w8(32'hbb963054),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c615e95),
	.w1(32'hbbcde7a8),
	.w2(32'hbbaee048),
	.w3(32'h3b8c800c),
	.w4(32'hbc81a067),
	.w5(32'h3d763174),
	.w6(32'h3b5c3df2),
	.w7(32'h38b176d8),
	.w8(32'h3d22f158),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f25455),
	.w1(32'h3b73f65d),
	.w2(32'h3b2d8d7a),
	.w3(32'hbc109d15),
	.w4(32'hbc38b022),
	.w5(32'h3abafa3c),
	.w6(32'hbc4221fc),
	.w7(32'h3c192fa4),
	.w8(32'hbbe73e41),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc03224a),
	.w1(32'h3d1d46a1),
	.w2(32'h3cf23ae8),
	.w3(32'h3b29e3dd),
	.w4(32'h38ef87eb),
	.w5(32'hba617d8d),
	.w6(32'hbb81523a),
	.w7(32'h3b983a63),
	.w8(32'h3c1afde5),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c13e9bd),
	.w1(32'h3bcab1ff),
	.w2(32'h3b3bf85a),
	.w3(32'h3ba37cae),
	.w4(32'hb953a2da),
	.w5(32'hbc0a9cc9),
	.w6(32'hbc95cd84),
	.w7(32'h3ca777e6),
	.w8(32'hbc372dae),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9689aa),
	.w1(32'h3cbadde7),
	.w2(32'h3b1072e7),
	.w3(32'hbc6541ee),
	.w4(32'h3d2257f4),
	.w5(32'hbc4db7d9),
	.w6(32'h3c54757e),
	.w7(32'hbb93e627),
	.w8(32'h3b38f61f),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7d4002),
	.w1(32'hbac67718),
	.w2(32'h3b5ed110),
	.w3(32'h3bfb1a75),
	.w4(32'hbc9ae0bf),
	.w5(32'hbbd4a4ec),
	.w6(32'hbb42c4d1),
	.w7(32'h3a675c3b),
	.w8(32'hbc08215e),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc374f7a),
	.w1(32'hbbdf5915),
	.w2(32'h3b76d77d),
	.w3(32'hbc618169),
	.w4(32'hb91de014),
	.w5(32'hbbc46e1a),
	.w6(32'h3b872a7b),
	.w7(32'hbc0d5057),
	.w8(32'hbbb6d465),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd06308a),
	.w1(32'hbc8c039b),
	.w2(32'h3c33492a),
	.w3(32'hbc223d64),
	.w4(32'hbc967160),
	.w5(32'hbc60cc12),
	.w6(32'hbbf808aa),
	.w7(32'h3b42c820),
	.w8(32'hba9d1a6f),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcebbc63),
	.w1(32'hbb7ef4d4),
	.w2(32'hbb661630),
	.w3(32'h3b9f0889),
	.w4(32'h3b87ad99),
	.w5(32'hba89e0c6),
	.w6(32'h3a9f2305),
	.w7(32'hbc0d0ea9),
	.w8(32'h3bd5358f),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c20c111),
	.w1(32'hbbd6ba91),
	.w2(32'hbb54c50f),
	.w3(32'h3d31b8a8),
	.w4(32'hb9a4ae4a),
	.w5(32'hbb3ebb96),
	.w6(32'h3be43201),
	.w7(32'h3b8dbdb2),
	.w8(32'hbcb9ba4d),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adc8e06),
	.w1(32'h3ca73d3a),
	.w2(32'hbc429fa1),
	.w3(32'h3bcaa98a),
	.w4(32'h3a762e6f),
	.w5(32'h3cf6a712),
	.w6(32'hba568234),
	.w7(32'hbb37fee7),
	.w8(32'hba730fdb),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4b5398),
	.w1(32'h3c8f5396),
	.w2(32'h3da06b6e),
	.w3(32'h3b97a827),
	.w4(32'h3c679af3),
	.w5(32'h3a07d7b5),
	.w6(32'h3abb260b),
	.w7(32'h3c8d3ba8),
	.w8(32'h3b3a1054),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3b0329),
	.w1(32'hbcdfb427),
	.w2(32'hbbca026e),
	.w3(32'hbb74f224),
	.w4(32'hbb1f2f0e),
	.w5(32'hbc0e55c5),
	.w6(32'hbb069138),
	.w7(32'hbca2c4ab),
	.w8(32'hbc01fc51),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b99fdde),
	.w1(32'hbabb1f91),
	.w2(32'hbba20ff1),
	.w3(32'h3c018ff2),
	.w4(32'hbbb74561),
	.w5(32'h3bd44ab7),
	.w6(32'hbc05bcca),
	.w7(32'h3b6d858c),
	.w8(32'h3aeb6b7a),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a99ea),
	.w1(32'hbc1a483d),
	.w2(32'h3b6fb729),
	.w3(32'hbc56ad79),
	.w4(32'h3c3bd9fc),
	.w5(32'h3c126c5a),
	.w6(32'h3cce52bb),
	.w7(32'hb99a7051),
	.w8(32'hbb253a08),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cf8ef2f),
	.w1(32'h3bc7a866),
	.w2(32'h3b2009a6),
	.w3(32'hbb321860),
	.w4(32'h3a469128),
	.w5(32'hba2c4dc9),
	.w6(32'hbc21fb7d),
	.w7(32'h3b6ca76b),
	.w8(32'h3bc604e6),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4a1ca6),
	.w1(32'h3afa8f95),
	.w2(32'hbc00ebed),
	.w3(32'hbbfe3b9c),
	.w4(32'h3b1b4499),
	.w5(32'hbce40a8b),
	.w6(32'hbb01965e),
	.w7(32'h3a938f4d),
	.w8(32'hbc8492d1),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4a4c6d),
	.w1(32'h3c0030a1),
	.w2(32'h3bd96af1),
	.w3(32'h3bd27e8d),
	.w4(32'hbc3a6f42),
	.w5(32'hbbb867f1),
	.w6(32'hbb035e46),
	.w7(32'hbc9546d0),
	.w8(32'h3b040659),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb46b9f),
	.w1(32'hbca98de0),
	.w2(32'hbb0ef3de),
	.w3(32'hba784c12),
	.w4(32'hbbff3df2),
	.w5(32'hbb015ab5),
	.w6(32'hbafec761),
	.w7(32'h38fa9785),
	.w8(32'hbccdcdb5),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba059a8),
	.w1(32'hbb871589),
	.w2(32'h3ca57740),
	.w3(32'hbc96b1ce),
	.w4(32'hba6ac7fa),
	.w5(32'hbbdb9264),
	.w6(32'hb9c26728),
	.w7(32'hbca1cc9f),
	.w8(32'h38949613),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0d59b9),
	.w1(32'h3cd6145d),
	.w2(32'hb9b2ed13),
	.w3(32'hbc524523),
	.w4(32'hbc2fb451),
	.w5(32'h3c1bcbe4),
	.w6(32'hbb8ecab0),
	.w7(32'hba5c87d1),
	.w8(32'h3a9874cf),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcde33ed),
	.w1(32'hbc817224),
	.w2(32'hbd0e1f92),
	.w3(32'h3b61b549),
	.w4(32'hbc38a8cc),
	.w5(32'hbcb53ef1),
	.w6(32'hb98513a6),
	.w7(32'h3c278a5b),
	.w8(32'h3b58c579),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdf8f2b),
	.w1(32'hbc071496),
	.w2(32'h3c1762ee),
	.w3(32'hba821e4e),
	.w4(32'hbc608d22),
	.w5(32'hbc921b6c),
	.w6(32'hbb66e313),
	.w7(32'hbad93561),
	.w8(32'hba272b10),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0e6b7c),
	.w1(32'hbbed4dc7),
	.w2(32'h3d062fa8),
	.w3(32'h3b6b67d5),
	.w4(32'h3b268d98),
	.w5(32'hbce57194),
	.w6(32'hbc31da37),
	.w7(32'h3c0e5e7c),
	.w8(32'hbc3b2ea4),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1d592a),
	.w1(32'hbb95891e),
	.w2(32'hbcb7cf30),
	.w3(32'h3bbed481),
	.w4(32'hbb8ace50),
	.w5(32'hbb567f87),
	.w6(32'hba137f89),
	.w7(32'hbbb6ec13),
	.w8(32'h3d48180b),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be197d0),
	.w1(32'h3b5f138a),
	.w2(32'hbc8eef44),
	.w3(32'hbbb55b76),
	.w4(32'hbc1c029b),
	.w5(32'hbc15b67f),
	.w6(32'hb9c3a2f1),
	.w7(32'hbbd6c03a),
	.w8(32'hbcd7c341),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc95ae69),
	.w1(32'h3b84a1cd),
	.w2(32'hbcd152da),
	.w3(32'hbc269963),
	.w4(32'hbc1d4198),
	.w5(32'h3c13a8eb),
	.w6(32'hbc196957),
	.w7(32'hbc2eff59),
	.w8(32'hbc86dcdf),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb06ce0),
	.w1(32'hba4ae61f),
	.w2(32'hbbf82430),
	.w3(32'h3b8df59c),
	.w4(32'h3be15ee6),
	.w5(32'hbb9f49da),
	.w6(32'h3b48dfcf),
	.w7(32'h3c2200e3),
	.w8(32'h3b11c6fc),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b375743),
	.w1(32'hbcf7d589),
	.w2(32'hbb483d63),
	.w3(32'hbbf1ebfa),
	.w4(32'h3c6dcc46),
	.w5(32'hbc8ff44c),
	.w6(32'h3c62eb45),
	.w7(32'h3c13c65d),
	.w8(32'h3bd65cb2),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc01425e),
	.w1(32'hbba45c2a),
	.w2(32'hbc815b3d),
	.w3(32'hbb2b031f),
	.w4(32'hbcbfc7d2),
	.w5(32'h3adf64c5),
	.w6(32'hbbf7fed3),
	.w7(32'h3baa0e4b),
	.w8(32'h3b8b5b83),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc155168),
	.w1(32'h3c2a48b8),
	.w2(32'hbc75fa41),
	.w3(32'h3d4e0244),
	.w4(32'h3c5b4c88),
	.w5(32'h3cec368e),
	.w6(32'hbbcc748b),
	.w7(32'hbc96b2e8),
	.w8(32'hbb8c6c19),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8c77da),
	.w1(32'hbc177211),
	.w2(32'hbb5efac7),
	.w3(32'hbcae8c9f),
	.w4(32'hbcad931c),
	.w5(32'h3baef6a9),
	.w6(32'hbb9ad2a2),
	.w7(32'h3c76000d),
	.w8(32'hbc06ea99),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9d0c64),
	.w1(32'hbb757298),
	.w2(32'hbb4cf769),
	.w3(32'hbbc7b363),
	.w4(32'h3b11fc08),
	.w5(32'hbc97eb93),
	.w6(32'hbc43a983),
	.w7(32'hbc522dc9),
	.w8(32'h3c03b1ca),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba8a9b2),
	.w1(32'hbc6b6c41),
	.w2(32'h3ba16050),
	.w3(32'hbc4e6660),
	.w4(32'h3b9ba04b),
	.w5(32'h3bbe8e35),
	.w6(32'hbc108bb9),
	.w7(32'hbbc9bd83),
	.w8(32'h3bd445d0),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394d4eb9),
	.w1(32'h3af1604a),
	.w2(32'hbd080cf9),
	.w3(32'hbb276769),
	.w4(32'hbcdd6803),
	.w5(32'hbcca5066),
	.w6(32'hbc229f55),
	.w7(32'hbc855b7f),
	.w8(32'hbc1fea4b),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0bbe0f),
	.w1(32'h3c246387),
	.w2(32'hbd23fcff),
	.w3(32'h3b91d3f3),
	.w4(32'hba7870ad),
	.w5(32'hbce4c081),
	.w6(32'h3c99417d),
	.w7(32'hbb6a710f),
	.w8(32'h3827dae4),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8f5d5b),
	.w1(32'h3b86b919),
	.w2(32'hbcd44b86),
	.w3(32'hbc8bbf0d),
	.w4(32'h3c4e2991),
	.w5(32'h3c5f2edd),
	.w6(32'hbb886d6f),
	.w7(32'h39e62638),
	.w8(32'h3b9d08f7),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb918d0d7),
	.w1(32'h3a8e8d64),
	.w2(32'h3c26760c),
	.w3(32'h3a8eb9a2),
	.w4(32'hbc887d5b),
	.w5(32'hbb900338),
	.w6(32'hbc32c883),
	.w7(32'hbc461c7e),
	.w8(32'hbbdce8a1),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4e58b9),
	.w1(32'h3aad8dcd),
	.w2(32'h3c244de7),
	.w3(32'h3c8192d8),
	.w4(32'h3b88533e),
	.w5(32'h3c124db1),
	.w6(32'h3b4db21a),
	.w7(32'hbcdccc7b),
	.w8(32'hba367d6e),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba11c704),
	.w1(32'hbbf5375a),
	.w2(32'h3c23b2d8),
	.w3(32'hbc80dc02),
	.w4(32'hbce0d472),
	.w5(32'hbc4b0b92),
	.w6(32'hbc1e97ce),
	.w7(32'hbb0a2123),
	.w8(32'h3c4a1243),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0ed4c2),
	.w1(32'h3b037bd3),
	.w2(32'hbc9f7641),
	.w3(32'h3d0fd79a),
	.w4(32'h39186f60),
	.w5(32'h3bce6eeb),
	.w6(32'h3b781fd8),
	.w7(32'h3bd80072),
	.w8(32'h3abf3fda),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8e77b5),
	.w1(32'h3b5223d8),
	.w2(32'h3bbb5d47),
	.w3(32'hb9ac7f0d),
	.w4(32'h3b525ed7),
	.w5(32'hbb08057a),
	.w6(32'hbc2e3061),
	.w7(32'hbbf4fbd9),
	.w8(32'hbc4f7216),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc80b801),
	.w1(32'h392e2791),
	.w2(32'h3cb90767),
	.w3(32'hbd20f2e9),
	.w4(32'h3c85cccc),
	.w5(32'hba77cf72),
	.w6(32'hb86041c1),
	.w7(32'h3a9b6132),
	.w8(32'h3c1d1017),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d9a93),
	.w1(32'hbb8d6495),
	.w2(32'hbabcdfc8),
	.w3(32'hbc7bccbb),
	.w4(32'h3d553937),
	.w5(32'h3cb4d947),
	.w6(32'h3a90d3b3),
	.w7(32'h3bbc3a95),
	.w8(32'h3a1cb086),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b435df4),
	.w1(32'h3c6030c0),
	.w2(32'hbbf7e480),
	.w3(32'h3b2d6e66),
	.w4(32'hbb6810f6),
	.w5(32'h39cf16e5),
	.w6(32'hbc1f83ed),
	.w7(32'hbbc5f720),
	.w8(32'hbc28c9b5),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1566fe),
	.w1(32'hbca06e0c),
	.w2(32'hbc3ca048),
	.w3(32'hbcf506a8),
	.w4(32'hbbcb42ec),
	.w5(32'h3c64b680),
	.w6(32'hbd107ea5),
	.w7(32'h3a4f67e5),
	.w8(32'hbc0cf2db),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf6153a),
	.w1(32'h3b8eb468),
	.w2(32'hbb7d1b28),
	.w3(32'hbbe477b0),
	.w4(32'hbc329e72),
	.w5(32'hbbd4a875),
	.w6(32'h3b7e4244),
	.w7(32'hba140ae0),
	.w8(32'hbbfb41cf),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1e8678),
	.w1(32'hbc3c55d9),
	.w2(32'hbc697fd8),
	.w3(32'hbbecf175),
	.w4(32'h3d180d0f),
	.w5(32'h3b713e35),
	.w6(32'hbb5d6818),
	.w7(32'hbad72e13),
	.w8(32'hbca58bf3),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc285653),
	.w1(32'h3bbefe72),
	.w2(32'hbc07933c),
	.w3(32'h3d25d3ba),
	.w4(32'h3c8bd80f),
	.w5(32'hbb03f506),
	.w6(32'hbc92894b),
	.w7(32'hbc3cef6f),
	.w8(32'hbb73e55d),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9dc79c),
	.w1(32'hba949a20),
	.w2(32'h3b56fa15),
	.w3(32'h3bf4408f),
	.w4(32'h3b9db5e4),
	.w5(32'hbb8a5129),
	.w6(32'h3a9cdd88),
	.w7(32'h3d0a5850),
	.w8(32'hbbdcf0a4),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1050fe),
	.w1(32'hbb060493),
	.w2(32'h3c75e33f),
	.w3(32'hbbb6d7cd),
	.w4(32'hbb519b13),
	.w5(32'hba4d5fef),
	.w6(32'hbbca705c),
	.w7(32'h3bc5378f),
	.w8(32'h3b4c387a),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba82e93),
	.w1(32'h3c0b21c3),
	.w2(32'hbc0ca6ef),
	.w3(32'hbbf5b5ae),
	.w4(32'hbc257de8),
	.w5(32'hbb6b6bc7),
	.w6(32'h3a229bd1),
	.w7(32'h3bad0550),
	.w8(32'h3b114634),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7994e6),
	.w1(32'hbb905680),
	.w2(32'hbb2aa1d7),
	.w3(32'h3cac7ce1),
	.w4(32'h3c5f5c8e),
	.w5(32'h3b1a1a4d),
	.w6(32'hbadc2969),
	.w7(32'hbb93c7d0),
	.w8(32'hbbd09796),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c16c2e2),
	.w1(32'hbadb52f1),
	.w2(32'hbbba9995),
	.w3(32'h3b8c1df9),
	.w4(32'h3a9e78e0),
	.w5(32'h3a776bcc),
	.w6(32'hba26b295),
	.w7(32'hbbc7fab6),
	.w8(32'h3b589fbf),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb096898),
	.w1(32'h3afd82bd),
	.w2(32'hbc4ab959),
	.w3(32'hbc0aaa4e),
	.w4(32'hba6bf56c),
	.w5(32'h39ccf206),
	.w6(32'h3cc617d7),
	.w7(32'hbb29ad88),
	.w8(32'hbbd7a375),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb824bd8),
	.w1(32'hbbe7d699),
	.w2(32'hba882140),
	.w3(32'h3adb8aff),
	.w4(32'h39cec25a),
	.w5(32'hbbbae293),
	.w6(32'hbbbadfbf),
	.w7(32'hbb1c90f7),
	.w8(32'hbbce1535),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a8e51),
	.w1(32'h39b01b39),
	.w2(32'h3b8a62bf),
	.w3(32'h3b5c7c75),
	.w4(32'hba0e4f99),
	.w5(32'h3b8d7def),
	.w6(32'hbb3eacc2),
	.w7(32'hbbd8e314),
	.w8(32'hbb997d85),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd07ab0d),
	.w1(32'hba425911),
	.w2(32'hbab0b6f4),
	.w3(32'h3b0e8e45),
	.w4(32'h3ad08f21),
	.w5(32'hbc382fda),
	.w6(32'h3b3e38cd),
	.w7(32'h3b3f5fa7),
	.w8(32'hbb464d19),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7a7aa0),
	.w1(32'h3d274e3c),
	.w2(32'hb80f68db),
	.w3(32'h3bdc33e4),
	.w4(32'h3bef6a49),
	.w5(32'h3b9c5b7b),
	.w6(32'hba8c086e),
	.w7(32'h3bc0a35e),
	.w8(32'hbbb3ac48),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbe969e),
	.w1(32'h3b7af19a),
	.w2(32'hba35b322),
	.w3(32'hbc0fa6b6),
	.w4(32'h3abf013d),
	.w5(32'hbade3e88),
	.w6(32'h3b43001d),
	.w7(32'h3c2ef1b0),
	.w8(32'h3b88d536),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b233b56),
	.w1(32'h3c12617d),
	.w2(32'hbbe08173),
	.w3(32'h3c863d74),
	.w4(32'h3c5f2e91),
	.w5(32'h3b1cf13f),
	.w6(32'hba22316f),
	.w7(32'h3c802bdc),
	.w8(32'h3c492ea3),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc58ea67),
	.w1(32'h3b44a713),
	.w2(32'h3b9545a5),
	.w3(32'h3be0aa07),
	.w4(32'h3b598a06),
	.w5(32'h3c50f6b7),
	.w6(32'h3d612038),
	.w7(32'hbc1baeaf),
	.w8(32'h3b417f7d),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bba83b5),
	.w1(32'hbc0573de),
	.w2(32'h3b3d9ac4),
	.w3(32'hbb4e1bae),
	.w4(32'hb9d1579e),
	.w5(32'h3b11f50f),
	.w6(32'h3b8545a6),
	.w7(32'h36def89d),
	.w8(32'hbbf44510),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb115c68),
	.w1(32'h3baff543),
	.w2(32'h3bcd0f5b),
	.w3(32'hbc5267ac),
	.w4(32'h3c4abed6),
	.w5(32'hbc201f3d),
	.w6(32'h3ba81e1e),
	.w7(32'hbbae9e34),
	.w8(32'h3c26eb0d),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7f77f8),
	.w1(32'hbb0c97e8),
	.w2(32'hbb59b352),
	.w3(32'h3d598dcb),
	.w4(32'hbb39fa71),
	.w5(32'hbc25fdb3),
	.w6(32'hbb4f132c),
	.w7(32'hbcb60008),
	.w8(32'hbc41286a),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7086a6),
	.w1(32'h3ac4b7ed),
	.w2(32'hbc28aa59),
	.w3(32'h3c0bcd37),
	.w4(32'hbba15bc1),
	.w5(32'hbb646588),
	.w6(32'hbbfef9d7),
	.w7(32'h3b8af085),
	.w8(32'hbc43b445),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2d69ae),
	.w1(32'hbb667a04),
	.w2(32'hbb06cbeb),
	.w3(32'hbabba45e),
	.w4(32'h398a92d5),
	.w5(32'h3cc01220),
	.w6(32'hbb05ffe7),
	.w7(32'hbbc1978b),
	.w8(32'h3a4855bc),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b08f364),
	.w1(32'hb96622c6),
	.w2(32'h3c8f8ffb),
	.w3(32'h3bd33a00),
	.w4(32'hbb610b55),
	.w5(32'hba93467d),
	.w6(32'hbc98c7b1),
	.w7(32'h3b00097d),
	.w8(32'h3bc8b13e),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc27dbfe),
	.w1(32'hbce40dd4),
	.w2(32'hbb9890b4),
	.w3(32'h3c72d4eb),
	.w4(32'hbcc8b2d2),
	.w5(32'hbc43fee4),
	.w6(32'h3cb07ab5),
	.w7(32'h3b8a9440),
	.w8(32'hba74da18),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc600b22),
	.w1(32'h3ac11132),
	.w2(32'h3be32948),
	.w3(32'hba1bfb31),
	.w4(32'hbc525078),
	.w5(32'hbb22078d),
	.w6(32'hbc7d3935),
	.w7(32'hbc0e78e8),
	.w8(32'hbc2327bf),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c86e7b2),
	.w1(32'hbbd29c60),
	.w2(32'hbb5d3f4d),
	.w3(32'h3c0dc49f),
	.w4(32'h3b83d661),
	.w5(32'hbbf231bd),
	.w6(32'hbbc34343),
	.w7(32'h3bd66390),
	.w8(32'h3c624fe2),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba71216),
	.w1(32'hbbdedba3),
	.w2(32'h3c3fa1bb),
	.w3(32'h3bac74fa),
	.w4(32'hbbf94e66),
	.w5(32'h3bb7ba65),
	.w6(32'hbb95d7cb),
	.w7(32'h3be3ac43),
	.w8(32'hbae45b41),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a08ce16),
	.w1(32'hba328591),
	.w2(32'hbc51962d),
	.w3(32'h3ca57dd3),
	.w4(32'hbae6c0da),
	.w5(32'h3b4930c6),
	.w6(32'hbc8bdf59),
	.w7(32'hbbcd1724),
	.w8(32'h3b5aa687),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b51bf80),
	.w1(32'hbb944182),
	.w2(32'hbb339ecb),
	.w3(32'h3bd260ef),
	.w4(32'hbb313f99),
	.w5(32'hbc23256e),
	.w6(32'h3ab4d526),
	.w7(32'h3c8434d5),
	.w8(32'hbb8a9c9f),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c93beb),
	.w1(32'hbb9bbd13),
	.w2(32'hbb790304),
	.w3(32'hbc613cdd),
	.w4(32'hbbd1333f),
	.w5(32'h3adc5d9e),
	.w6(32'hbb9818f5),
	.w7(32'hbad1e88d),
	.w8(32'hbb1b100b),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2336a4),
	.w1(32'hbcc7fbff),
	.w2(32'h3a50a9b7),
	.w3(32'h3a19e09e),
	.w4(32'h3c13a43f),
	.w5(32'hbcf9a313),
	.w6(32'hbbd274a0),
	.w7(32'hbc113b1c),
	.w8(32'hbb2067c5),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbb2ff0),
	.w1(32'hbad45256),
	.w2(32'hb8917991),
	.w3(32'h3b3a0ac1),
	.w4(32'hbc8eea6e),
	.w5(32'hbc5e3333),
	.w6(32'h3b403451),
	.w7(32'h3c885edb),
	.w8(32'hbc0f773e),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc40cc6),
	.w1(32'h3b32c037),
	.w2(32'hbebed6e7),
	.w3(32'hba082d88),
	.w4(32'h3bbd3f44),
	.w5(32'hbef39299),
	.w6(32'hbc6b8ef0),
	.w7(32'hbf1fedde),
	.w8(32'hbf4265bb),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ee781fe),
	.w1(32'hbf15d721),
	.w2(32'hbf8aff3a),
	.w3(32'hbf1a2a5a),
	.w4(32'h3b8f4dd8),
	.w5(32'hbf066e55),
	.w6(32'hbf395c01),
	.w7(32'hbf09d33b),
	.w8(32'hbf3420da),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbf45db06),
	.w1(32'hbee772a5),
	.w2(32'hbf0b0822),
	.w3(32'hbf381651),
	.w4(32'hbf072da2),
	.w5(32'hbf05ed26),
	.w6(32'hbf135f0b),
	.w7(32'hbe268761),
	.w8(32'hbf0073ce),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbef1e46b),
	.w1(32'hbe9dc41d),
	.w2(32'hbf1f48fc),
	.w3(32'hbe8e8a83),
	.w4(32'hbf2e37d5),
	.w5(32'hbea7e9b0),
	.w6(32'hbee763b7),
	.w7(32'hbf167087),
	.w8(32'hbf3143a2),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbf2a2aff),
	.w1(32'hbf168932),
	.w2(32'hbf3ce20d),
	.w3(32'hbf1921b9),
	.w4(32'hbe99f816),
	.w5(32'hbf3fffb4),
	.w6(32'hbef71cf6),
	.w7(32'hbf8dc9f1),
	.w8(32'hbeef69f5),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9ad84c),
	.w1(32'hbf9d2ba2),
	.w2(32'hbe628ff7),
	.w3(32'hbf1be453),
	.w4(32'hbf38c938),
	.w5(32'hbf0fb767),
	.w6(32'hbf054e35),
	.w7(32'hbf573156),
	.w8(32'hbf2988fb),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbead86f6),
	.w1(32'hbec873b4),
	.w2(32'hbf8794db),
	.w3(32'hbee90a6c),
	.w4(32'hbf3a0ece),
	.w5(32'hbe9af87b),
	.w6(32'hbef484fc),
	.w7(32'hbf149575),
	.w8(32'hbf04e62c),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbf1cf53e),
	.w1(32'hbf08d1b5),
	.w2(32'hbf3a0509),
	.w3(32'hbf099fef),
	.w4(32'hbeb0185a),
	.w5(32'hbf1024e0),
	.w6(32'hbf86c93c),
	.w7(32'hbee047ed),
	.w8(32'hbf28dace),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbf4c44c4),
	.w1(32'hbf10d72e),
	.w2(32'hbe907824),
	.w3(32'hbf08974e),
	.w4(32'hbf158bf9),
	.w5(32'hbf81f0bd),
	.w6(32'hbe5f401a),
	.w7(32'hbf19d195),
	.w8(32'hbf0054fa),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbf15452a),
	.w1(32'hbee1adbc),
	.w2(32'hbeda5bd9),
	.w3(32'hbec34c0c),
	.w4(32'hbf1a063f),
	.w5(32'hbf169769),
	.w6(32'hbf4cd00e),
	.w7(32'hbf0135d8),
	.w8(32'hbec0c8de),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbe5d66dd),
	.w1(32'h3dcc4d30),
	.w2(32'hbf72b6c8),
	.w3(32'hbf5645ab),
	.w4(32'hbf47166e),
	.w5(32'hbf1367c0),
	.w6(32'hbec25e64),
	.w7(32'hbeef00a4),
	.w8(32'hbf0cfc3e),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbe94601f),
	.w1(32'hbf8444e9),
	.w2(32'hbf3517bb),
	.w3(32'hbf3adf96),
	.w4(32'hbf02ea76),
	.w5(32'hbf45a21b),
	.w6(32'hbe82ad34),
	.w7(32'hbee117e2),
	.w8(32'hbe1bba0e),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbf844bef),
	.w1(32'hbf0c2d48),
	.w2(32'hbef6954d),
	.w3(32'hbee60f94),
	.w4(32'hbf07ae6f),
	.w5(32'hbe336fec),
	.w6(32'hbf0a4ee7),
	.w7(32'hbf1f36ec),
	.w8(32'hbeea2854),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbf0066ff),
	.w1(32'hbfb79d66),
	.w2(32'hbf20622b),
	.w3(32'hbf87f75d),
	.w4(32'hbf12b7bc),
	.w5(32'hbf2897a2),
	.w6(32'hbef7e04b),
	.w7(32'hbebd175c),
	.w8(32'hbf0da0e3),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbf951f78),
	.w1(32'hbf6ed506),
	.w2(32'hbf0502c4),
	.w3(32'hbebae298),
	.w4(32'hbef69f76),
	.w5(32'hbf057086),
	.w6(32'hbf5fb985),
	.w7(32'hbee89d0a),
	.w8(32'hbec326e1),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbf02e11b),
	.w1(32'hbed06fd9),
	.w2(32'hbec87ed6),
	.w3(32'hbf373175),
	.w4(32'hbec17f24),
	.w5(32'hbf50e30d),
	.w6(32'hbf297ae5),
	.w7(32'hbf70d909),
	.w8(32'hbf2d57cb),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbf258ad5),
	.w1(32'hbf119562),
	.w2(32'hbef0d7b8),
	.w3(32'hbf24c05f),
	.w4(32'hbf235315),
	.w5(32'hbed864b3),
	.w6(32'hbf16a80c),
	.w7(32'hbeef038a),
	.w8(32'hbf87c371),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbf304ef9),
	.w1(32'hbf3cf8e2),
	.w2(32'hbf10a12e),
	.w3(32'hbee1d1b0),
	.w4(32'hbfaf3715),
	.w5(32'hbea35f79),
	.w6(32'hbef95522),
	.w7(32'hbf7fed1c),
	.w8(32'hbf412822),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbf0e11b0),
	.w1(32'hbf840a1e),
	.w2(32'hbeef7baa),
	.w3(32'hbf1ed98c),
	.w4(32'hbf2c1bfe),
	.w5(32'hbf215cfd),
	.w6(32'hbf05ef34),
	.w7(32'hbf3ab99a),
	.w8(32'hbed1888f),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbf05afce),
	.w1(32'hbdc829e1),
	.w2(32'hbf04efd2),
	.w3(32'hbec33b16),
	.w4(32'hbf188de5),
	.w5(32'h3eeb1af7),
	.w6(32'hbf1d553b),
	.w7(32'hbf08d3a9),
	.w8(32'hbf6648c6),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbf361b70),
	.w1(32'hbf056394),
	.w2(32'hbf3c2712),
	.w3(32'hbf024700),
	.w4(32'hbee283c3),
	.w5(32'hbf4bb9da),
	.w6(32'hbf4f7992),
	.w7(32'hbf387930),
	.w8(32'hbf086ded),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbeb7567a),
	.w1(32'hbed3c8cb),
	.w2(32'hbf4afb29),
	.w3(32'hbf4aa3f7),
	.w4(32'hbf13b5ab),
	.w5(32'hbed3c790),
	.w6(32'hbf0be89f),
	.w7(32'hbf1f665e),
	.w8(32'hbf0a7123),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbf07e3b4),
	.w1(32'hbefdf2f1),
	.w2(32'hbeb6bce4),
	.w3(32'hbee775a2),
	.w4(32'hbe47794c),
	.w5(32'hbf142ca0),
	.w6(32'hbef5678c),
	.w7(32'hbf29c1ad),
	.w8(32'hbf5819aa),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbf6187cb),
	.w1(32'hbedaeaa2),
	.w2(32'hbf7aad49),
	.w3(32'hbf12e07e),
	.w4(32'hbf12c1fb),
	.w5(32'hbed21f9e),
	.w6(32'hbefedb37),
	.w7(32'hbe476517),
	.w8(32'hbe6ae8c4),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbf11bea9),
	.w1(32'hbf1e6b62),
	.w2(32'hbe8cde3b),
	.w3(32'hbec4c9d2),
	.w4(32'hbeb022fd),
	.w5(32'hbf3fda7f),
	.w6(32'hbf1b4370),
	.w7(32'hbf03f897),
	.w8(32'hbeda9a30),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbf3b7b44),
	.w1(32'hbf5e11a0),
	.w2(32'hbef2b2cc),
	.w3(32'hbf52c3e4),
	.w4(32'hbe8b3caa),
	.w5(32'hbf1ff9a8),
	.w6(32'hbee270a4),
	.w7(32'hbf03598c),
	.w8(32'hbf23362a),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbf1530eb),
	.w1(32'hbefd55ad),
	.w2(32'hbf3031b2),
	.w3(32'hbedce451),
	.w4(32'hbe62eeb8),
	.w5(32'hbf4218e2),
	.w6(32'hbf1a6335),
	.w7(32'hbe266b31),
	.w8(32'hbf13635a),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbe971806),
	.w1(32'hbecca4c6),
	.w2(32'hbeabf4f7),
	.w3(32'hbf296028),
	.w4(32'hbedfe6b4),
	.w5(32'hbf1d4812),
	.w6(32'hbed721f3),
	.w7(32'hbe22bacd),
	.w8(32'hbf0646d3),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbe71c82b),
	.w1(32'hbf05cb4a),
	.w2(32'hbeccca9f),
	.w3(32'hbeeb3339),
	.w4(32'hbf4472ed),
	.w5(32'hbedfee99),
	.w6(32'hbf1a0ea9),
	.w7(32'hbed1badc),
	.w8(32'hbf0ca913),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f65c5ca),
	.w1(32'h3dcdefea),
	.w2(32'h3f48059a),
	.w3(32'h3f7328ff),
	.w4(32'h3f96df24),
	.w5(32'h37f0edbc),
	.w6(32'h36a1459d),
	.w7(32'h37031aaa),
	.w8(32'h3e9f4e93),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f1abf3c),
	.w1(32'h3d372030),
	.w2(32'hb6eb99d8),
	.w3(32'h3f56cd17),
	.w4(32'h3fa2eaf0),
	.w5(32'h3efbfd2f),
	.w6(32'h3f04dc08),
	.w7(32'h3ee12fdb),
	.w8(32'h3f87f5e2),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f2bcdc4),
	.w1(32'h3f26d6ee),
	.w2(32'h3e2c3e79),
	.w3(32'h38a4e302),
	.w4(32'h3f5a6ba4),
	.w5(32'h3f34b648),
	.w6(32'h3ec7709e),
	.w7(32'h3e8c043e),
	.w8(32'h368e8a83),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f2c38d5),
	.w1(32'h3f00ddd6),
	.w2(32'h3dcc240e),
	.w3(32'h3f0557b0),
	.w4(32'h3fb746c2),
	.w5(32'h3f0cf8a4),
	.w6(32'h3df1b6bf),
	.w7(32'h3edfca97),
	.w8(32'h3f02cba8),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f883e69),
	.w1(32'h3f24f1ea),
	.w2(32'h3f1934c1),
	.w3(32'h3e9d6ebe),
	.w4(32'h3ef15464),
	.w5(32'h3f81c582),
	.w6(32'h3efc3932),
	.w7(32'hb72eb61b),
	.w8(32'h3f4e357c),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f4397af),
	.w1(32'h3ebd1ac9),
	.w2(32'hb7adc04e),
	.w3(32'h3eda33a6),
	.w4(32'h33bffb8f),
	.w5(32'h3ebb7ca5),
	.w6(32'h3f35b3af),
	.w7(32'h3f2f817a),
	.w8(32'h3fafee1a),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f3b75f2),
	.w1(32'h391737a9),
	.w2(32'h3f85650c),
	.w3(32'h3f86071d),
	.w4(32'h34193b06),
	.w5(32'h3eedc7e4),
	.w6(32'h3ee40df9),
	.w7(32'h389da508),
	.w8(32'h3cb39543),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3e86a202),
	.w1(32'h3f44b783),
	.w2(32'h3ee25338),
	.w3(32'h3f96b2a5),
	.w4(32'h3ee26d8c),
	.w5(32'h3f9de5b1),
	.w6(32'h3f9074f0),
	.w7(32'h3ec0219b),
	.w8(32'h3f4e1bd7),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f2aff81),
	.w1(32'h363b73a8),
	.w2(32'h3efffafa),
	.w3(32'h36ab4346),
	.w4(32'h3f27c921),
	.w5(32'hb73577d2),
	.w6(32'h3f9e3e13),
	.w7(32'h3ee33ac6),
	.w8(32'h3f033b95),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ecc4b76),
	.w1(32'h3f09dc1e),
	.w2(32'h3eff0b9f),
	.w3(32'h3e818dc6),
	.w4(32'h3f1953f8),
	.w5(32'h3ed699b9),
	.w6(32'h3f138fbf),
	.w7(32'h35a70a87),
	.w8(32'h3d65075d),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f260790),
	.w1(32'h3ec4f25b),
	.w2(32'h3f588cbb),
	.w3(32'h3fd4da7f),
	.w4(32'h3ed4a510),
	.w5(32'h3f75dc72),
	.w6(32'h3d06e252),
	.w7(32'h3ef0ff2a),
	.w8(32'h3c9844ea),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f884f5c),
	.w1(32'h3eb074e6),
	.w2(32'hb6afc828),
	.w3(32'h3fa36de9),
	.w4(32'h3f6a4caf),
	.w5(32'h3eb91296),
	.w6(32'h3f3e942f),
	.w7(32'h3eca6c83),
	.w8(32'h37789502),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f0c16c2),
	.w1(32'h3ea645e5),
	.w2(32'h3eac96f3),
	.w3(32'h3f27ae4d),
	.w4(32'h3e88db9c),
	.w5(32'h3ffcccb1),
	.w6(32'h3ebdcdc8),
	.w7(32'h3f844826),
	.w8(32'h3ef5d022),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d57eb6f),
	.w1(32'h3d09eff8),
	.w2(32'h3f3770d9),
	.w3(32'h330dc92e),
	.w4(32'h3f901bda),
	.w5(32'h3f4a74f2),
	.w6(32'h3f9c96f9),
	.w7(32'h3de32abe),
	.w8(32'h3eb92a6a),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3e95c708),
	.w1(32'h3ec433e8),
	.w2(32'h3f949b4c),
	.w3(32'h3da9921d),
	.w4(32'h3ee9fff1),
	.w5(32'h3f5691fd),
	.w6(32'h3e2520b4),
	.w7(32'h3f79a3ce),
	.w8(32'h3ec1883d),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f718c6a),
	.w1(32'h3fc12320),
	.w2(32'h3f03aaf2),
	.w3(32'h3f29be72),
	.w4(32'h3f343978),
	.w5(32'h3f8f43f9),
	.w6(32'h3f9bb9b9),
	.w7(32'h3f664975),
	.w8(32'h36e302b2),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ed4fbea),
	.w1(32'h3d407fe2),
	.w2(32'h3f8ece1a),
	.w3(32'h3ea9618d),
	.w4(32'h3bc6bbb7),
	.w5(32'h3efee8da),
	.w6(32'h3f1ff997),
	.w7(32'hb7be69ca),
	.w8(32'h3fd0214c),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f3a8f16),
	.w1(32'h3f3b8755),
	.w2(32'h3f41e181),
	.w3(32'h3e8288e7),
	.w4(32'h3e78af90),
	.w5(32'h3f0b27b4),
	.w6(32'h3ea4a160),
	.w7(32'h3e0b61eb),
	.w8(32'h3f071c3f),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f0c4947),
	.w1(32'h3ec0e998),
	.w2(32'h33a6957d),
	.w3(32'h3e9dcb13),
	.w4(32'h3c41e352),
	.w5(32'h3ed2af2e),
	.w6(32'hb595eb3c),
	.w7(32'h3f81e6e2),
	.w8(32'h3efda13a),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3edda313),
	.w1(32'h3f7158ad),
	.w2(32'h3e9de179),
	.w3(32'h3f4ed447),
	.w4(32'h3f03d3ec),
	.w5(32'h3e28fa87),
	.w6(32'h3f79b820),
	.w7(32'h3e520f0d),
	.w8(32'h3f002ee1),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3e93da77),
	.w1(32'h3f8b8316),
	.w2(32'hb5dd57fc),
	.w3(32'h3f08c1c2),
	.w4(32'h3f0b51e6),
	.w5(32'h3f07c930),
	.w6(32'h3e1c2447),
	.w7(32'h3f6a0aa3),
	.w8(32'h3fa666f8),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3eea0368),
	.w1(32'h3d4c9d56),
	.w2(32'h3f24a1e3),
	.w3(32'h3f49095c),
	.w4(32'h3edf6c21),
	.w5(32'h3e81dda3),
	.w6(32'h3f3375f4),
	.w7(32'h3e80e715),
	.w8(32'hb5562805),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f660fb0),
	.w1(32'h3f34313c),
	.w2(32'h3f004c20),
	.w3(32'h3e1c933e),
	.w4(32'h3f61ba2e),
	.w5(32'h3eb92f5c),
	.w6(32'h36b1af23),
	.w7(32'h3e96019e),
	.w8(32'h3e2b963b),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f414576),
	.w1(32'h3dc9d0a2),
	.w2(32'h3e3c1b35),
	.w3(32'h3f692143),
	.w4(32'h3e9e32b9),
	.w5(32'h3f2bd1dc),
	.w6(32'h3ec693a0),
	.w7(32'h3f044713),
	.w8(32'hb5babf13),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3e2f2249),
	.w1(32'h3eaaa6b7),
	.w2(32'h3f2dfdf4),
	.w3(32'h3f5a9caf),
	.w4(32'h3f932755),
	.w5(32'h3f9acabc),
	.w6(32'h3eb9109b),
	.w7(32'h3f16e0f4),
	.w8(32'h3ec3e0cb),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3e81ba20),
	.w1(32'h3f8fe1bf),
	.w2(32'h3df8a48e),
	.w3(32'h3ec184e0),
	.w4(32'h3f1d273d),
	.w5(32'h3ead338c),
	.w6(32'h3f0af41d),
	.w7(32'h3e5e6dc4),
	.w8(32'h3d139194),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6ee9385),
	.w1(32'h3bed193c),
	.w2(32'h3f97cb31),
	.w3(32'h3f4df76a),
	.w4(32'h3e953214),
	.w5(32'h3ed2ba61),
	.w6(32'h3f725618),
	.w7(32'h3f3f1fae),
	.w8(32'h3f22b13e),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3f2c1175),
	.w1(32'h3ef6b372),
	.w2(32'h3ee3ce40),
	.w3(32'h3e76291a),
	.w4(32'h3ed5190f),
	.w5(32'h3e08f937),
	.w6(32'h3ee0cd8d),
	.w7(32'hb65c2eaa),
	.w8(32'h3f0970fa),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca75d0e),
	.w1(32'h3f0abbe2),
	.w2(32'hb60753d2),
	.w3(32'h3f98807f),
	.w4(32'h3df081cd),
	.w5(32'h3d124fd7),
	.w6(32'h351ec30d),
	.w7(32'h3d426623),
	.w8(32'h3ce46536),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3601409f),
	.w1(32'h3cdb3817),
	.w2(32'hbdacd1a8),
	.w3(32'hbce3e89c),
	.w4(32'hbd3ef94c),
	.w5(32'h3cb167c5),
	.w6(32'hb8aa198c),
	.w7(32'h3b4c3e20),
	.w8(32'hbc0b2f94),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d675c20),
	.w1(32'h3d72e77e),
	.w2(32'h3d064e29),
	.w3(32'hb612b14b),
	.w4(32'h3d762d65),
	.w5(32'h3de7038b),
	.w6(32'h3cec895a),
	.w7(32'h368c7f98),
	.w8(32'h3d38db1b),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbe701fac),
	.w1(32'h361fd14e),
	.w2(32'h3d48d60b),
	.w3(32'h3cb88e4f),
	.w4(32'h3dc04cec),
	.w5(32'h3e06cbce),
	.w6(32'h3dda87ba),
	.w7(32'h3e1ad6b5),
	.w8(32'hbcad14fa),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd01503e),
	.w1(32'hbd0e8e89),
	.w2(32'hbeb6e259),
	.w3(32'h3c7d3765),
	.w4(32'h3e100a43),
	.w5(32'h3cd5a1ee),
	.w6(32'h3c25b68e),
	.w7(32'h3d983304),
	.w8(32'h3cc5573d),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97bf092),
	.w1(32'hbd9c0789),
	.w2(32'h3d144c08),
	.w3(32'h3d2e08fb),
	.w4(32'h3d88b2fd),
	.w5(32'hbce53ac5),
	.w6(32'h3d8b6c43),
	.w7(32'h3d208272),
	.w8(32'hb6a34606),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbb357b),
	.w1(32'h3dc6ac6e),
	.w2(32'hbda790cd),
	.w3(32'h3935a677),
	.w4(32'h3c572255),
	.w5(32'h394fd952),
	.w6(32'hbb86a4aa),
	.w7(32'h3af5c4e2),
	.w8(32'hb682036b),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38aab517),
	.w1(32'h3c87b2f9),
	.w2(32'h3d473760),
	.w3(32'h3dee63be),
	.w4(32'h3d30995d),
	.w5(32'h3d95c002),
	.w6(32'h3a94eeda),
	.w7(32'hbd16771d),
	.w8(32'h3d732416),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbe42264d),
	.w1(32'hbcde3f6a),
	.w2(32'h3ce6ad9d),
	.w3(32'h3daee86e),
	.w4(32'h3d36505c),
	.w5(32'hb89694ba),
	.w6(32'h3b67a818),
	.w7(32'h38aaae82),
	.w8(32'hbcc45b68),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3e1fca72),
	.w1(32'h3ca29504),
	.w2(32'h3cf28949),
	.w3(32'hbdce0fac),
	.w4(32'h3ddc6624),
	.w5(32'hbdd03606),
	.w6(32'hb75031d8),
	.w7(32'h3b73d77e),
	.w8(32'hbcc37969),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb75c90c3),
	.w1(32'h3c11317e),
	.w2(32'h3cf9a706),
	.w3(32'h3e1b9cbd),
	.w4(32'hbd9fb486),
	.w5(32'h3db15c02),
	.w6(32'hbc090c97),
	.w7(32'h3d8df860),
	.w8(32'h3d9c2356),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d7eaed6),
	.w1(32'hbc0b9839),
	.w2(32'h3cb9b6e5),
	.w3(32'hbe31926d),
	.w4(32'h3dab29ec),
	.w5(32'h3c9f791f),
	.w6(32'h3d9c5ea7),
	.w7(32'h3dae4f8b),
	.w8(32'hbce4b364),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cec7cf4),
	.w1(32'hb846b1fb),
	.w2(32'hbccab084),
	.w3(32'h38515fb0),
	.w4(32'hbd9d5e5b),
	.w5(32'h3cb8eab2),
	.w6(32'h3d3fc203),
	.w7(32'h3da6e5d0),
	.w8(32'hbc200fee),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d92d9af),
	.w1(32'hbbaf35b3),
	.w2(32'h3dd63ca7),
	.w3(32'h3dec814c),
	.w4(32'h3b139f21),
	.w5(32'h3c4c2a39),
	.w6(32'h3d2085a6),
	.w7(32'hb61479e1),
	.w8(32'h3e48c575),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf7496b),
	.w1(32'h3bc575b3),
	.w2(32'h3d2532e7),
	.w3(32'h399f2882),
	.w4(32'hba93d1b6),
	.w5(32'h3cf82489),
	.w6(32'hbc6596f1),
	.w7(32'h3d17503c),
	.w8(32'h3d058434),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3f98a7),
	.w1(32'h3d672061),
	.w2(32'h3b4d7e5d),
	.w3(32'h3d976eed),
	.w4(32'hbdb52ffa),
	.w5(32'hbe0aaa19),
	.w6(32'h3ca9450d),
	.w7(32'hbda1f64b),
	.w8(32'h3da42607),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb84c573),
	.w1(32'hb7bb9564),
	.w2(32'hb9e8aa04),
	.w3(32'h3ce146c0),
	.w4(32'hbcfc89c7),
	.w5(32'h3d198b52),
	.w6(32'h3d08291d),
	.w7(32'hbbbee3e7),
	.w8(32'h3bb06a5d),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7764e6f),
	.w1(32'hbdb3074f),
	.w2(32'h3d48a26f),
	.w3(32'hbcd1676e),
	.w4(32'hbc12e2fe),
	.w5(32'hbd0cde2b),
	.w6(32'h3d398cde),
	.w7(32'hbbd90551),
	.w8(32'h3d9216cf),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cf6076b),
	.w1(32'hbd8bde49),
	.w2(32'hb4425937),
	.w3(32'hbd3d4e17),
	.w4(32'h3cb9049b),
	.w5(32'h3d98d4f8),
	.w6(32'h3dff4cc4),
	.w7(32'h3d0f6689),
	.w8(32'h3c8dc1f7),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbdbd601a),
	.w1(32'h3d4b82d8),
	.w2(32'h3e0326c6),
	.w3(32'h35aeff5d),
	.w4(32'h3c78d1cb),
	.w5(32'h3df932f4),
	.w6(32'hbd077099),
	.w7(32'h3d828d09),
	.w8(32'hbcf62431),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cf19a24),
	.w1(32'h3cd3810c),
	.w2(32'h3d17cb19),
	.w3(32'h3d3f5322),
	.w4(32'h3d45667a),
	.w5(32'h3d2ed21e),
	.w6(32'h3bb0fa4c),
	.w7(32'hbe6dc1cf),
	.w8(32'h3cd0b706),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbe1f33d8),
	.w1(32'h3c8e65ec),
	.w2(32'h3d07614a),
	.w3(32'h35fa7153),
	.w4(32'h3c27d89e),
	.w5(32'hbabf6cbf),
	.w6(32'h3e228afb),
	.w7(32'h3d9f5435),
	.w8(32'h3de78f32),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b88d0cb),
	.w1(32'hb5a80cbd),
	.w2(32'hb57563e5),
	.w3(32'h3d90cbf9),
	.w4(32'hbe224c34),
	.w5(32'h3dd26f0f),
	.w6(32'h3cdfff3c),
	.w7(32'h3d0247cc),
	.w8(32'h3e5186b8),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbd4b7f),
	.w1(32'h3d2402e0),
	.w2(32'hbd073e57),
	.w3(32'h3d8d1ec2),
	.w4(32'h3e107160),
	.w5(32'h3d3ce7ce),
	.w6(32'hbd9836bc),
	.w7(32'h3d39bd02),
	.w8(32'h3c8b2669),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbdd6c6ad),
	.w1(32'h34bceca8),
	.w2(32'h3d4cc7ea),
	.w3(32'h3d20dc43),
	.w4(32'h3d64c8d5),
	.w5(32'hbb54a33e),
	.w6(32'h3ca11b2a),
	.w7(32'hbda7e8cd),
	.w8(32'h3d94c95d),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbe470c1f),
	.w1(32'h3de2039e),
	.w2(32'h3b3d0827),
	.w3(32'hbcde66d6),
	.w4(32'hbd233594),
	.w5(32'h3c986cf4),
	.w6(32'hbcd9e3f7),
	.w7(32'h3dab5423),
	.w8(32'hbc5b4aa7),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d8b0045),
	.w1(32'h3c155bc5),
	.w2(32'hbcb4e522),
	.w3(32'h3d000c0c),
	.w4(32'h35c3d7cf),
	.w5(32'h39e58b6f),
	.w6(32'hbd154ab4),
	.w7(32'h3dd79cd0),
	.w8(32'hbbeb811a),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cebe667),
	.w1(32'h3dac504f),
	.w2(32'h3dafafcb),
	.w3(32'h3ceb66a0),
	.w4(32'h3d03aebd),
	.w5(32'hbd19ebfc),
	.w6(32'h3c9a7b47),
	.w7(32'h3d39d613),
	.w8(32'hbd16e01b),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6012698),
	.w1(32'h3c87faa4),
	.w2(32'hb71e9b88),
	.w3(32'h3d05e84b),
	.w4(32'h3c3ad49f),
	.w5(32'h3d0d8073),
	.w6(32'h3d7eadf6),
	.w7(32'h3dc99def),
	.w8(32'h3d0e1471),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d1f69a6),
	.w1(32'h3dcb5dca),
	.w2(32'h35f01ff6),
	.w3(32'h34c2d684),
	.w4(32'h3588c870),
	.w5(32'h3d464403),
	.w6(32'h3ab6c45e),
	.w7(32'h3ccf7478),
	.w8(32'h3d1617f3),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c149083),
	.w1(32'h3d42d4c3),
	.w2(32'h3c75f0e7),
	.w3(32'h3c53cbe3),
	.w4(32'h3c090d85),
	.w5(32'h3d22c3a2),
	.w6(32'h39ede32c),
	.w7(32'hb620bf22),
	.w8(32'h3d168fde),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3585baee),
	.w1(32'h3d013629),
	.w2(32'h3ca26700),
	.w3(32'h3c326f8c),
	.w4(32'h3d107f0c),
	.w5(32'h35632d9e),
	.w6(32'h3cb15485),
	.w7(32'h3aec503a),
	.w8(32'h3c8efc5f),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5fd9f4),
	.w1(32'h3db220de),
	.w2(32'h3c7d1b45),
	.w3(32'h3abf85a9),
	.w4(32'h3c1fdb56),
	.w5(32'h3cb411dc),
	.w6(32'h3c7a69a2),
	.w7(32'h3a86d67d),
	.w8(32'h3d0c4554),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b69b730),
	.w1(32'h3d06977c),
	.w2(32'h3cf8acfd),
	.w3(32'h3c53c542),
	.w4(32'h32d44ece),
	.w5(32'h3d2cf3d8),
	.w6(32'h3cb657fe),
	.w7(32'h3c52a0f7),
	.w8(32'h3cdb4c93),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d0cbb00),
	.w1(32'hb6745633),
	.w2(32'h3c24a0c2),
	.w3(32'h3d0ee28e),
	.w4(32'h3cc40692),
	.w5(32'h3d72798a),
	.w6(32'h3bf1e943),
	.w7(32'hb69d4d95),
	.w8(32'h3c9e4d4c),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce0fcf6),
	.w1(32'hb2ed6e84),
	.w2(32'h3c3efda3),
	.w3(32'h3c5c8232),
	.w4(32'h334b00b6),
	.w5(32'h3949cd36),
	.w6(32'h344aefc2),
	.w7(32'h3d3d2f1b),
	.w8(32'h3c5a632f),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d826904),
	.w1(32'h3c05dd6f),
	.w2(32'h3d392ee8),
	.w3(32'h3d23967c),
	.w4(32'h3c0e4730),
	.w5(32'h3d15f46e),
	.w6(32'h3cc3a69f),
	.w7(32'h3cb0082b),
	.w8(32'h3cc19c92),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h33605eb2),
	.w1(32'h3c9d4cd3),
	.w2(32'hb1be744c),
	.w3(32'h3d185cb8),
	.w4(32'h3c2a32da),
	.w5(32'h3c5b55df),
	.w6(32'h3405f68d),
	.w7(32'h3c91dfe8),
	.w8(32'h3c117bb9),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bacad0d),
	.w1(32'h3cb5138b),
	.w2(32'h3ce430a3),
	.w3(32'h3c7dab4f),
	.w4(32'hb3f8893b),
	.w5(32'h3a309f81),
	.w6(32'h3cb930bc),
	.w7(32'h3c92c2ea),
	.w8(32'h3cb7e5d4),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d94406d),
	.w1(32'h3cb7d48d),
	.w2(32'h3cf6ef6a),
	.w3(32'h3a0b69dc),
	.w4(32'h3c0ff0c1),
	.w5(32'h38a72ef0),
	.w6(32'h3be577ce),
	.w7(32'h3d2addb7),
	.w8(32'h3d503d37),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d235ce4),
	.w1(32'h3d096f38),
	.w2(32'h3c337711),
	.w3(32'h3cd8bd85),
	.w4(32'h3c03f412),
	.w5(32'hb5c03d36),
	.w6(32'h3ca441b0),
	.w7(32'hb357cc3a),
	.w8(32'h3c6ce0cb),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbd25d7),
	.w1(32'h3b8d31bb),
	.w2(32'h3da7cffb),
	.w3(32'h3d060c7c),
	.w4(32'h3c727511),
	.w5(32'h3c60e6c9),
	.w6(32'h3b9f05fa),
	.w7(32'h3bd4f423),
	.w8(32'h3a3dc7a5),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb2d57349),
	.w1(32'h3d164974),
	.w2(32'h3cc3dfe1),
	.w3(32'h3d3b68bf),
	.w4(32'h3a442447),
	.w5(32'h3c1bd92e),
	.w6(32'h39aef419),
	.w7(32'h3cb519cd),
	.w8(32'h3bcb6426),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a53c58c),
	.w1(32'h3c3099fc),
	.w2(32'h3ca5fa66),
	.w3(32'h3b056c9a),
	.w4(32'h3d567976),
	.w5(32'h3c46d4d9),
	.w6(32'h3c991461),
	.w7(32'h3d54ec3e),
	.w8(32'h3d354880),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9a2df7),
	.w1(32'h3d07271e),
	.w2(32'h3db06772),
	.w3(32'h3d2ad36d),
	.w4(32'h3cfe0dab),
	.w5(32'h351ffcf8),
	.w6(32'h3db55c71),
	.w7(32'h3c827225),
	.w8(32'h3c50abf1),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd23e07),
	.w1(32'h38207545),
	.w2(32'h3c1994d6),
	.w3(32'h3cac8d2d),
	.w4(32'h34ae05bb),
	.w5(32'h3d7618e2),
	.w6(32'h3a51b56b),
	.w7(32'h3d5b1dac),
	.w8(32'h3c864a7f),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b78f219),
	.w1(32'h3b2b163a),
	.w2(32'h3be9a61f),
	.w3(32'h3be4a829),
	.w4(32'h3b11866d),
	.w5(32'h3c53847c),
	.w6(32'h3cbf2fc1),
	.w7(32'h3cc7422f),
	.w8(32'h3c43e53e),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0e9a25),
	.w1(32'h39506e87),
	.w2(32'h3c8bfc8f),
	.w3(32'hb53ee891),
	.w4(32'h3d7c7860),
	.w5(32'h3c495c4e),
	.w6(32'h3c18032d),
	.w7(32'hb5989bc2),
	.w8(32'h3c66d173),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cafcc6d),
	.w1(32'h3c85c9d7),
	.w2(32'h3b05f676),
	.w3(32'h3d9ecd5a),
	.w4(32'h3b33399b),
	.w5(32'h3c8f6e9c),
	.w6(32'h3d22bc57),
	.w7(32'h3b3d8921),
	.w8(32'h3bd45ce3),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d10f9b7),
	.w1(32'h3c8417b0),
	.w2(32'h3c2570c2),
	.w3(32'h3ae57739),
	.w4(32'h3d5c19bb),
	.w5(32'h3d7ffacc),
	.w6(32'h3d846e4f),
	.w7(32'h3377aafa),
	.w8(32'h3c296c14),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cae31ec),
	.w1(32'h3c3abd53),
	.w2(32'h3b92e8ac),
	.w3(32'h3cf9a830),
	.w4(32'h3ba6b381),
	.w5(32'h33b4ecd8),
	.w6(32'h39eb7ac6),
	.w7(32'h3cc1c8df),
	.w8(32'h3d834765),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aadc235),
	.w1(32'h3cd8277d),
	.w2(32'h3c49ccd8),
	.w3(32'h32af6d3b),
	.w4(32'h3b9114ac),
	.w5(32'h3b138bb9),
	.w6(32'h3cb84bbf),
	.w7(32'h3c6ad539),
	.w8(32'h3d74b99c),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d0b13b9),
	.w1(32'h3b9c6603),
	.w2(32'h3ca4f7e4),
	.w3(32'h3c1a8710),
	.w4(32'h3c9045e0),
	.w5(32'h328e4517),
	.w6(32'h3aee95a8),
	.w7(32'h3aab8c30),
	.w8(32'h3b136eb4),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d2e944c),
	.w1(32'h3d3004c9),
	.w2(32'h3d596640),
	.w3(32'h3baf79d5),
	.w4(32'h3ca4936e),
	.w5(32'h3c72ee3e),
	.w6(32'h3c01ade8),
	.w7(32'h3cc83cfc),
	.w8(32'h3b7d4690),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2d1021),
	.w1(32'h3c992f4a),
	.w2(32'h3bca0e11),
	.w3(32'h3c3583be),
	.w4(32'h3b1f127a),
	.w5(32'h3a05c856),
	.w6(32'h3d982461),
	.w7(32'h3a925078),
	.w8(32'hb67a729a),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d10e9dc),
	.w1(32'h3c16647f),
	.w2(32'h3c7ced13),
	.w3(32'h3d491ab5),
	.w4(32'h3cbcf3f6),
	.w5(32'h3cd3ad23),
	.w6(32'h384d5103),
	.w7(32'h3da3c742),
	.w8(32'h3d4f6b64),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b91cdd8),
	.w1(32'h3c8cebf1),
	.w2(32'h3ae25b40),
	.w3(32'h3cadc8d2),
	.w4(32'h3608dcd4),
	.w5(32'h3c5abd70),
	.w6(32'h3c09c09a),
	.w7(32'h3c1978e1),
	.w8(32'h397b85e1),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d97c3d8),
	.w1(32'hbb3601b8),
	.w2(32'hbb56d369),
	.w3(32'hb5cdbb9b),
	.w4(32'hbc523457),
	.w5(32'hbc8836b0),
	.w6(32'h3ca0db9f),
	.w7(32'hbbcbc7a7),
	.w8(32'hbbb58ca1),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdcb69f),
	.w1(32'hbb4d932b),
	.w2(32'hbb68abf2),
	.w3(32'hbb9b73ea),
	.w4(32'hbbbf3a55),
	.w5(32'hbbff84ca),
	.w6(32'hbbfb8230),
	.w7(32'hbb970e04),
	.w8(32'h3c604840),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb48ef2f),
	.w1(32'hbb551f1b),
	.w2(32'hbc122505),
	.w3(32'hbc01d70c),
	.w4(32'h3bac0d60),
	.w5(32'h3cdac34b),
	.w6(32'h3bd879a4),
	.w7(32'hb8b8ba7b),
	.w8(32'hbc5be5ba),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb62f247),
	.w1(32'hbb891594),
	.w2(32'hbb753b2b),
	.w3(32'hbb4f04d1),
	.w4(32'hbc75f9f7),
	.w5(32'hbbd918a2),
	.w6(32'hbc376693),
	.w7(32'hbbd25182),
	.w8(32'hbbde304f),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8f501b),
	.w1(32'hbad41081),
	.w2(32'h3a9ab889),
	.w3(32'hbc11fc00),
	.w4(32'hba83e6d7),
	.w5(32'h3a8fff7e),
	.w6(32'hbbb31175),
	.w7(32'h3b6deb04),
	.w8(32'hbbc1e3b8),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8e943c),
	.w1(32'hbc976527),
	.w2(32'hbc79e203),
	.w3(32'hbb57e5ae),
	.w4(32'hbc843cef),
	.w5(32'hbc3f1779),
	.w6(32'h3a63291f),
	.w7(32'hbc8a02a6),
	.w8(32'hbc8c35c9),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc13c64a),
	.w1(32'h3bfb8367),
	.w2(32'h3bdae2ce),
	.w3(32'hbc9fc236),
	.w4(32'h3c46bb8e),
	.w5(32'h3c526951),
	.w6(32'hbba4cb5d),
	.w7(32'hbab9209a),
	.w8(32'hbb66c84c),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2186ca),
	.w1(32'h3b83d199),
	.w2(32'h3c2da1f7),
	.w3(32'hb994fe01),
	.w4(32'h3c005fab),
	.w5(32'hbad1c107),
	.w6(32'h3b1a8d4c),
	.w7(32'h3c087d56),
	.w8(32'h3a119da9),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b923a34),
	.w1(32'hbc1ebf82),
	.w2(32'hbc494986),
	.w3(32'h3c2f7866),
	.w4(32'hbb25803d),
	.w5(32'h3cd1bbd5),
	.w6(32'hb8505a41),
	.w7(32'h3baa78db),
	.w8(32'h3b0a51e9),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa085f6),
	.w1(32'h3b20f577),
	.w2(32'h3c0556bd),
	.w3(32'h3a1d0cfa),
	.w4(32'h3aa377e9),
	.w5(32'h3b9090d6),
	.w6(32'h3b4fd1b5),
	.w7(32'h397d1e65),
	.w8(32'hbb8baa7d),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0b8be2),
	.w1(32'h3bc8a460),
	.w2(32'h3c0350f0),
	.w3(32'h3b957a3f),
	.w4(32'hbbd45951),
	.w5(32'hbc64b1ca),
	.w6(32'h3ac0b4a8),
	.w7(32'h3c11d79a),
	.w8(32'h3c123f5b),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37b6fb3c),
	.w1(32'h3bf95f51),
	.w2(32'h3c2004ac),
	.w3(32'h3b833111),
	.w4(32'hbbad3756),
	.w5(32'hbc240d44),
	.w6(32'hbb091c4b),
	.w7(32'h3b762430),
	.w8(32'hbab5f1ab),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8a5d53),
	.w1(32'h3c044045),
	.w2(32'h3b5017af),
	.w3(32'hbb06ff75),
	.w4(32'h3a86d5d3),
	.w5(32'hba8a7d73),
	.w6(32'hbb06bb88),
	.w7(32'h3a645e9e),
	.w8(32'h3b283033),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba825416),
	.w1(32'h3b38b20f),
	.w2(32'h3aab8624),
	.w3(32'h3b3457c9),
	.w4(32'h3be91a74),
	.w5(32'h3b3c658a),
	.w6(32'h3ab545ca),
	.w7(32'h3b92a7d2),
	.w8(32'h3c21e7f3),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b216099),
	.w1(32'hbab78995),
	.w2(32'h3bfddd93),
	.w3(32'h3a934788),
	.w4(32'hbc6e711e),
	.w5(32'hbcc256e7),
	.w6(32'h3bfa7924),
	.w7(32'h39943499),
	.w8(32'h3c282a02),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb0b893),
	.w1(32'h3b4bddd5),
	.w2(32'h3a412ded),
	.w3(32'hbc230f9b),
	.w4(32'h3b18c244),
	.w5(32'h3c92aa47),
	.w6(32'h3c3cf0ec),
	.w7(32'hbc346c08),
	.w8(32'hbbba7d0e),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b24e39e),
	.w1(32'hbb6a9408),
	.w2(32'h3ae52410),
	.w3(32'h3b650c7e),
	.w4(32'hbb5e6938),
	.w5(32'hbc1478c5),
	.w6(32'h3abebcdc),
	.w7(32'hbc021e6d),
	.w8(32'hbc3bc77b),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac78253),
	.w1(32'h3bba3876),
	.w2(32'h3c4b7247),
	.w3(32'hba53fbb5),
	.w4(32'h3ab317c5),
	.w5(32'hb83b85cf),
	.w6(32'hbb5ed144),
	.w7(32'h3c1f240e),
	.w8(32'h3c39a013),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcb10b6),
	.w1(32'h3bc32251),
	.w2(32'h3c862e69),
	.w3(32'h3c97e7a6),
	.w4(32'hbb3b68da),
	.w5(32'h39ad0cb1),
	.w6(32'hb9a1e3fa),
	.w7(32'hba5e92a1),
	.w8(32'h3b71ac8b),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdd365b),
	.w1(32'hbb684092),
	.w2(32'h3bcfd4eb),
	.w3(32'hbb09d975),
	.w4(32'h3af056b1),
	.w5(32'h3a8d3ce7),
	.w6(32'hba12b9b4),
	.w7(32'h3b861d9d),
	.w8(32'h3b4cc5d5),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbedbed8),
	.w1(32'hbbcfa20c),
	.w2(32'h3b894c48),
	.w3(32'h3bb6dbbb),
	.w4(32'hbae260db),
	.w5(32'hbc049a15),
	.w6(32'h3beb302f),
	.w7(32'hbac11393),
	.w8(32'h3c221bbe),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6ec5d8),
	.w1(32'h3b02a6d1),
	.w2(32'hbba1bbd3),
	.w3(32'hbb1e4d60),
	.w4(32'hbbe7f6d2),
	.w5(32'hbbccb911),
	.w6(32'h3b710e09),
	.w7(32'hbbd19ac6),
	.w8(32'hbb59faa2),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeedaaa),
	.w1(32'h39735fb4),
	.w2(32'h3c6b533d),
	.w3(32'h38c4ae95),
	.w4(32'hbbe9344a),
	.w5(32'hbc473d50),
	.w6(32'h3bbde508),
	.w7(32'hbb8e9487),
	.w8(32'h3b506ba2),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb846500a),
	.w1(32'h3bc25164),
	.w2(32'h3c11000d),
	.w3(32'hbc02aded),
	.w4(32'h3b4ebfea),
	.w5(32'h3b420bc3),
	.w6(32'hbaa7ed59),
	.w7(32'hbb9a8c80),
	.w8(32'hb9922a72),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd04065),
	.w1(32'h3bfc3d41),
	.w2(32'h3c48b7b2),
	.w3(32'h3aa5bd24),
	.w4(32'hbad9b109),
	.w5(32'hba080dc5),
	.w6(32'hbb998620),
	.w7(32'h3bd9b8a0),
	.w8(32'h3c32f9aa),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c16e6db),
	.w1(32'hbc336c52),
	.w2(32'hba92b5ec),
	.w3(32'h3c6e2d8d),
	.w4(32'hbc1af26f),
	.w5(32'hbbe756a9),
	.w6(32'h3c288bf8),
	.w7(32'h3ad568c8),
	.w8(32'h3be215bc),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc35ec78),
	.w1(32'hbb84194b),
	.w2(32'hbb139685),
	.w3(32'hbbf76e5c),
	.w4(32'hbb6bb5ee),
	.w5(32'hb99379dc),
	.w6(32'hba845a5c),
	.w7(32'h3b134cb2),
	.w8(32'hbc09ddc2),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b027835),
	.w1(32'hba1a13ab),
	.w2(32'h37a915ad),
	.w3(32'h39a03cc9),
	.w4(32'hbb2d2203),
	.w5(32'h3a1bec45),
	.w6(32'h3b0db414),
	.w7(32'hbb7aab4d),
	.w8(32'hbab2a08c),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b37b67e),
	.w1(32'hbbe5ec93),
	.w2(32'hbbf700b4),
	.w3(32'hbab7eee5),
	.w4(32'hbb828317),
	.w5(32'hbc64bdf5),
	.w6(32'hbb83c529),
	.w7(32'hbb966b16),
	.w8(32'hbb36c299),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8d7c98),
	.w1(32'hba023f3e),
	.w2(32'hbb9797ab),
	.w3(32'hbb55821d),
	.w4(32'hbc309858),
	.w5(32'hbc2bdff9),
	.w6(32'hbbfec5f1),
	.w7(32'hbbf6cf7a),
	.w8(32'hbc026788),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc24beee),
	.w1(32'h3872facc),
	.w2(32'hbbbb41da),
	.w3(32'hbbad0191),
	.w4(32'h3d0823ad),
	.w5(32'h3d5720f0),
	.w6(32'hbc3194cd),
	.w7(32'h3a8e8cde),
	.w8(32'h3ba8917d),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aca1bf2),
	.w1(32'h3b1c5042),
	.w2(32'h3c1f9428),
	.w3(32'h3c8b09af),
	.w4(32'hbb640af5),
	.w5(32'hbb05b3d4),
	.w6(32'h3cab3763),
	.w7(32'h3b90655b),
	.w8(32'h3bba7f38),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b22b9b8),
	.w1(32'hbbd8dd6a),
	.w2(32'h3a0fa930),
	.w3(32'h3b731c4d),
	.w4(32'hbafbf631),
	.w5(32'h39c3f4ea),
	.w6(32'h3ae77b20),
	.w7(32'h3a6177ad),
	.w8(32'h3b5e23ef),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3f4fc7),
	.w1(32'hb804a71c),
	.w2(32'hbbab5589),
	.w3(32'h3b155ed8),
	.w4(32'hbbb3c7bb),
	.w5(32'h3b1dd885),
	.w6(32'h3b831223),
	.w7(32'hbb9284fc),
	.w8(32'hbb8abe00),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8524e1),
	.w1(32'hbb1b02fd),
	.w2(32'hbbc11ef0),
	.w3(32'hba55a8d1),
	.w4(32'h3af42704),
	.w5(32'h3b40f18e),
	.w6(32'hbb90cedb),
	.w7(32'h3a6b7823),
	.w8(32'h3a975892),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38fada88),
	.w1(32'h39a3ba0c),
	.w2(32'h3c400f2a),
	.w3(32'hbc19042b),
	.w4(32'hbc089607),
	.w5(32'hbb628874),
	.w6(32'hbb21c7a1),
	.w7(32'h3afd5819),
	.w8(32'hbb8a3e1a),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c05a9c7),
	.w1(32'h3b87332f),
	.w2(32'hb8e5505e),
	.w3(32'hbb1e1fb2),
	.w4(32'hbb027ed3),
	.w5(32'h3ab2326c),
	.w6(32'hbb125a01),
	.w7(32'h3ba6ca95),
	.w8(32'h3b847362),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b02faa4),
	.w1(32'h3ae0c914),
	.w2(32'hbac3d33d),
	.w3(32'h3c1b3ca7),
	.w4(32'h3b6ac4ca),
	.w5(32'hbb2ad9a2),
	.w6(32'h3b330a9e),
	.w7(32'hba164e9a),
	.w8(32'h3bb24d76),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9fa113),
	.w1(32'hbb888663),
	.w2(32'hbb66ae3e),
	.w3(32'h3a1a41eb),
	.w4(32'hbaf7d92c),
	.w5(32'hba97aef6),
	.w6(32'h3bcc3e2d),
	.w7(32'hbb72c9ae),
	.w8(32'hbbce1a3a),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39155e13),
	.w1(32'hb98267b7),
	.w2(32'hbac5f424),
	.w3(32'hbbfd7726),
	.w4(32'hbb51f589),
	.w5(32'hbb716ef1),
	.w6(32'hbc716764),
	.w7(32'h3b9d6f31),
	.w8(32'h3bf4051c),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac0e178),
	.w1(32'hb9d7a631),
	.w2(32'h3bfeea2b),
	.w3(32'hbb399294),
	.w4(32'hba604ae3),
	.w5(32'h3b829794),
	.w6(32'h3b3b85d8),
	.w7(32'h3b77773d),
	.w8(32'h3ad3ac7e),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9edb9f),
	.w1(32'h3b930f6b),
	.w2(32'h3a37cc19),
	.w3(32'h3b17d889),
	.w4(32'hbc3c1435),
	.w5(32'hbc27f82f),
	.w6(32'hba18b174),
	.w7(32'hbc48e836),
	.w8(32'hbc00eb30),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8d9881),
	.w1(32'hbb9af61d),
	.w2(32'h3a26f638),
	.w3(32'hbc37c953),
	.w4(32'h3a3dac50),
	.w5(32'hbbfe22b4),
	.w6(32'hbc057288),
	.w7(32'h3c14c5f6),
	.w8(32'hbb27bb51),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfd6edd),
	.w1(32'hbb7be386),
	.w2(32'hbc1386e4),
	.w3(32'h3b8ff81d),
	.w4(32'h3aede6e8),
	.w5(32'h3b0e07be),
	.w6(32'hbb1768de),
	.w7(32'hbb02aa44),
	.w8(32'hbc2f5100),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba03eaf),
	.w1(32'hbbbd6228),
	.w2(32'h3bdb238c),
	.w3(32'h389f9558),
	.w4(32'hbbd5c6e0),
	.w5(32'hbc74433d),
	.w6(32'hbab4da65),
	.w7(32'h3b839a3f),
	.w8(32'h3bbee5eb),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9f6536),
	.w1(32'hbb1513ae),
	.w2(32'h3b3e1ee2),
	.w3(32'hbb5454e2),
	.w4(32'hbb1db0ba),
	.w5(32'hbbd4e489),
	.w6(32'h3bd4044d),
	.w7(32'hbb8682c0),
	.w8(32'hbbc642fb),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab085ee),
	.w1(32'h3ae0981a),
	.w2(32'hbb0f5718),
	.w3(32'hbb131dfe),
	.w4(32'hba63d8cd),
	.w5(32'h38396b6d),
	.w6(32'hb9c37c4e),
	.w7(32'h3bdbea6c),
	.w8(32'h3aa1816b),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b954999),
	.w1(32'h3b5feeac),
	.w2(32'h381bf9c0),
	.w3(32'hb983890e),
	.w4(32'h3c20caea),
	.w5(32'h3bc6c047),
	.w6(32'h3a8e524d),
	.w7(32'h3ba6dffd),
	.w8(32'h3baac16e),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af45be3),
	.w1(32'h3a9e7326),
	.w2(32'hbc17c19c),
	.w3(32'h3c6d77fd),
	.w4(32'h3b735efe),
	.w5(32'h3bf17c28),
	.w6(32'h3c49b27b),
	.w7(32'hbabef094),
	.w8(32'hbb547b1c),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3c4b08),
	.w1(32'hbb1dd1da),
	.w2(32'hbb745936),
	.w3(32'h3c2196c0),
	.w4(32'hbc938db2),
	.w5(32'h3b5cf914),
	.w6(32'h3b73c7a0),
	.w7(32'hbbbec48e),
	.w8(32'hbc2738a9),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabbf240),
	.w1(32'hba66daa2),
	.w2(32'hbc02c7b9),
	.w3(32'hbc146a99),
	.w4(32'hbbaac00b),
	.w5(32'hbba231e1),
	.w6(32'hba91cee1),
	.w7(32'h3b401c91),
	.w8(32'hbaea1d75),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a167096),
	.w1(32'h3b81c7a4),
	.w2(32'h3c3001f5),
	.w3(32'h39d776e4),
	.w4(32'hbaf907d5),
	.w5(32'hbbc93059),
	.w6(32'hba5defc8),
	.w7(32'hbabad382),
	.w8(32'hbbbf3a6f),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba19bc25),
	.w1(32'hbb5d42b9),
	.w2(32'hb9a933a0),
	.w3(32'h3c005b7c),
	.w4(32'hbb5ca5b5),
	.w5(32'hbc83d777),
	.w6(32'h3b810516),
	.w7(32'h3c73964e),
	.w8(32'h3cef144e),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb51aeb4),
	.w1(32'h3ba31dca),
	.w2(32'h3c2dac88),
	.w3(32'h3c48c90e),
	.w4(32'hbb2d0db4),
	.w5(32'hbbb98896),
	.w6(32'h3bc3d372),
	.w7(32'hbaa8d8ce),
	.w8(32'h3b57e2e3),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba946dba),
	.w1(32'hbbf6127a),
	.w2(32'h3b12af50),
	.w3(32'hbb92ea8d),
	.w4(32'h3bf979bf),
	.w5(32'h3b052838),
	.w6(32'h3b856f57),
	.w7(32'h3ba156e8),
	.w8(32'h3b5f9be3),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaed5186),
	.w1(32'hbc3e8283),
	.w2(32'hbc2b78e5),
	.w3(32'h3b4e15b8),
	.w4(32'h3bc83e3c),
	.w5(32'h3cb3f37d),
	.w6(32'hbac75247),
	.w7(32'h3a06c081),
	.w8(32'hbb4f6691),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc455ced),
	.w1(32'hba0e0685),
	.w2(32'h3b126864),
	.w3(32'hbbceadc6),
	.w4(32'hbc1e478b),
	.w5(32'hbb42e6d8),
	.w6(32'h389781d8),
	.w7(32'hbc2fad16),
	.w8(32'hbbd030ba),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4906b2),
	.w1(32'hbc03c6f2),
	.w2(32'hbbccefd1),
	.w3(32'hbba990d8),
	.w4(32'h3b833667),
	.w5(32'h3becb8ce),
	.w6(32'hbb049306),
	.w7(32'hbc3c042c),
	.w8(32'hbbc45c9c),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcd6715),
	.w1(32'hbbc0fc24),
	.w2(32'h3b1383be),
	.w3(32'h3b2b6ab7),
	.w4(32'hbb91adf7),
	.w5(32'hbb656bd0),
	.w6(32'hbb925a8d),
	.w7(32'hbbd3ca95),
	.w8(32'hbbf80b77),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule