module layer_10_featuremap_374(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb909644),
	.w1(32'hbbadba53),
	.w2(32'hbc16744a),
	.w3(32'h3bd0b010),
	.w4(32'h399accbb),
	.w5(32'h3c01c2d1),
	.w6(32'hbc1ba974),
	.w7(32'h3cbee7e8),
	.w8(32'h39688080),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba35d9f),
	.w1(32'h3b52207c),
	.w2(32'h3ba7ae85),
	.w3(32'h3b42ca9a),
	.w4(32'h3b52454c),
	.w5(32'h39a626f3),
	.w6(32'hbbdff1ba),
	.w7(32'hbd27d2eb),
	.w8(32'h3b600d03),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce66858),
	.w1(32'hbabc7b19),
	.w2(32'h3c8d1235),
	.w3(32'h3c87e759),
	.w4(32'hbc9b02f4),
	.w5(32'h3c8996a7),
	.w6(32'hbc06ad03),
	.w7(32'hbb9c6b2a),
	.w8(32'h3ae2b202),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbfc30c),
	.w1(32'hbb7c7e4c),
	.w2(32'hbc1c9b1c),
	.w3(32'h3bc8e5a4),
	.w4(32'h3c15c043),
	.w5(32'h3a9aec4f),
	.w6(32'h3ca89d5d),
	.w7(32'h3baa5055),
	.w8(32'hbb06f392),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab1b234),
	.w1(32'hba50c753),
	.w2(32'hbb6cdd3d),
	.w3(32'h3a71eaf5),
	.w4(32'hbac82bc5),
	.w5(32'hb991be3a),
	.w6(32'h3bee7491),
	.w7(32'h3b90364d),
	.w8(32'h3bcef46c),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d056b98),
	.w1(32'h3a008f91),
	.w2(32'h3b8b2dae),
	.w3(32'h3be365e9),
	.w4(32'h3ba4487f),
	.w5(32'h3cc47fd9),
	.w6(32'hbb9786e8),
	.w7(32'hbbd01d16),
	.w8(32'h3c0e3164),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc31176a),
	.w1(32'hbbbb53c0),
	.w2(32'hbb567e24),
	.w3(32'hbd0bc6cc),
	.w4(32'hbc933abf),
	.w5(32'hbb833993),
	.w6(32'hbca1601e),
	.w7(32'h3ba9f017),
	.w8(32'h3b48b93d),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c972152),
	.w1(32'hbc0e608e),
	.w2(32'h3a8f8220),
	.w3(32'hbaed7f16),
	.w4(32'hbc2b3ccc),
	.w5(32'hbc10c0a1),
	.w6(32'h3b49e1fc),
	.w7(32'h3c3a497a),
	.w8(32'hbc4dadf5),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3b8c60),
	.w1(32'h3bad7c0b),
	.w2(32'hbc18593b),
	.w3(32'h3c465e1d),
	.w4(32'hbc03476b),
	.w5(32'h3be6ae47),
	.w6(32'hbc1671be),
	.w7(32'hbaf6b63e),
	.w8(32'h3b23bb9f),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc567386),
	.w1(32'hba19b282),
	.w2(32'hbbfcfa12),
	.w3(32'hbbf047b6),
	.w4(32'hbbcf71d0),
	.w5(32'hbbad21d6),
	.w6(32'hbc567aeb),
	.w7(32'hbc14ffe1),
	.w8(32'h393a0e80),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb63194d),
	.w1(32'h3c01bda9),
	.w2(32'h3afdb051),
	.w3(32'h3c850dea),
	.w4(32'h3b7dc4af),
	.w5(32'hb9b9d9ba),
	.w6(32'h3afaf455),
	.w7(32'h3b856399),
	.w8(32'hbb835c8a),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c018b66),
	.w1(32'h3b88b2fa),
	.w2(32'h3b686a1c),
	.w3(32'h3c5925ac),
	.w4(32'hbd125ba3),
	.w5(32'hb99924f4),
	.w6(32'h3c32c8fa),
	.w7(32'h3b2eeaf1),
	.w8(32'h3c21ea3c),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb15c80),
	.w1(32'h3bb17a49),
	.w2(32'hbc1fc5e1),
	.w3(32'h3c36ab2d),
	.w4(32'hbbc75648),
	.w5(32'hbce3ed53),
	.w6(32'h3c2851e8),
	.w7(32'h3a39d558),
	.w8(32'h3b0e4d00),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1250b5),
	.w1(32'h3c4a9d32),
	.w2(32'h3c8603e3),
	.w3(32'hbc346db3),
	.w4(32'hbbaf55ce),
	.w5(32'h3af2844a),
	.w6(32'hbbb2a39f),
	.w7(32'h3ae55d3c),
	.w8(32'hbbc33d50),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8677dd),
	.w1(32'hba204b1c),
	.w2(32'hba4f00b3),
	.w3(32'hbce1ac28),
	.w4(32'hbbcaa851),
	.w5(32'h3c8f1f9c),
	.w6(32'hbc20340d),
	.w7(32'hbb9661de),
	.w8(32'h3a8cbdcd),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbca1f84),
	.w1(32'hbb15e97b),
	.w2(32'hbc058d35),
	.w3(32'h3b88f8c7),
	.w4(32'hb96ed2b5),
	.w5(32'h3a82b89d),
	.w6(32'hbc8460fb),
	.w7(32'h3bdd4cb8),
	.w8(32'hbb362510),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4d9d86),
	.w1(32'h3bf455ff),
	.w2(32'h3ba61bc2),
	.w3(32'hbb71c5bf),
	.w4(32'h3987ed54),
	.w5(32'hbbc4298d),
	.w6(32'hbb500437),
	.w7(32'h3b98ed77),
	.w8(32'h3bf78356),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaff8955),
	.w1(32'hbc21f32f),
	.w2(32'hbc5f4a54),
	.w3(32'hbcb3a4f3),
	.w4(32'hbc6ced2a),
	.w5(32'h3bfc14e3),
	.w6(32'h3d15362f),
	.w7(32'h3bc1e7f6),
	.w8(32'h3c1d69f5),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9abc85),
	.w1(32'hbc502874),
	.w2(32'hbc0ea888),
	.w3(32'h3c7f01e2),
	.w4(32'hbc5658e6),
	.w5(32'hbcd4fe4d),
	.w6(32'h3a9d8d2d),
	.w7(32'h3c303b34),
	.w8(32'h3b8b707d),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc4b5c9),
	.w1(32'hbb95c99d),
	.w2(32'h38c11bfc),
	.w3(32'hbc03df1b),
	.w4(32'hbab35aff),
	.w5(32'h3c973194),
	.w6(32'hbbd666c3),
	.w7(32'hbc76fbea),
	.w8(32'hbc4a1da8),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bacf3bc),
	.w1(32'h3a962211),
	.w2(32'h3c21f16c),
	.w3(32'hbc818cba),
	.w4(32'hbc5b23fc),
	.w5(32'hbb7e8e2d),
	.w6(32'h3a4e5b19),
	.w7(32'hbb5f542d),
	.w8(32'hbc879a32),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc11a47a),
	.w1(32'h3c907fc8),
	.w2(32'hbb8b2345),
	.w3(32'h3b6133fb),
	.w4(32'h3b912863),
	.w5(32'hbbc2e110),
	.w6(32'hbba86e5c),
	.w7(32'hbaba9901),
	.w8(32'hbc539135),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cfedd3b),
	.w1(32'hbc2feae9),
	.w2(32'hbc8f2753),
	.w3(32'h3b12196c),
	.w4(32'hbab9ae1d),
	.w5(32'h3b440463),
	.w6(32'h3a66ea95),
	.w7(32'h3ca6b3df),
	.w8(32'h3cd05e6e),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5cbda7),
	.w1(32'h399305c6),
	.w2(32'h3ca2bd4d),
	.w3(32'hbbc19c89),
	.w4(32'hbc004ae7),
	.w5(32'h39eae016),
	.w6(32'hbb53f17a),
	.w7(32'h398a91d1),
	.w8(32'h3ca4b8a6),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6d4a07),
	.w1(32'h3c36e58d),
	.w2(32'h3cbf6b0a),
	.w3(32'hbc044666),
	.w4(32'hbc38e962),
	.w5(32'h3b95dc8a),
	.w6(32'hbc0beb6d),
	.w7(32'h3c275b91),
	.w8(32'hbc78c1bc),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc84b084),
	.w1(32'hbb126c08),
	.w2(32'h3c855324),
	.w3(32'hbc0f0e77),
	.w4(32'hbbdb23b4),
	.w5(32'hbba82c48),
	.w6(32'h3b5b182e),
	.w7(32'h3b03b65e),
	.w8(32'hbc07af3b),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9acafbe),
	.w1(32'h38953657),
	.w2(32'h3beb236c),
	.w3(32'hbbd16fcd),
	.w4(32'h3cbc5b2b),
	.w5(32'hbc284390),
	.w6(32'h3abede65),
	.w7(32'hbb275308),
	.w8(32'h3bc0059e),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7e40c9),
	.w1(32'h3bb84755),
	.w2(32'hbb95f5b4),
	.w3(32'h3c2ba7b2),
	.w4(32'h3c0f95e3),
	.w5(32'hbdbffbe4),
	.w6(32'hbca11c2d),
	.w7(32'hbc660f24),
	.w8(32'hbc1a2432),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb299761),
	.w1(32'hbaa23deb),
	.w2(32'h3c32959d),
	.w3(32'hbad1b584),
	.w4(32'h3b731ecc),
	.w5(32'hbb40c908),
	.w6(32'h3baaa1ab),
	.w7(32'h3a174748),
	.w8(32'h3b3667d5),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ee3597),
	.w1(32'h3c70591c),
	.w2(32'h3c0277cd),
	.w3(32'hbb1bbc78),
	.w4(32'h3c9aad18),
	.w5(32'hbb108c75),
	.w6(32'hbc5432fa),
	.w7(32'hbc8aa734),
	.w8(32'hbba319f3),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5d9fcb),
	.w1(32'h3b876ab1),
	.w2(32'hbc1fae01),
	.w3(32'hbd69e063),
	.w4(32'hba9b5b99),
	.w5(32'h3b6de350),
	.w6(32'h3bdc4c69),
	.w7(32'hbb1417f9),
	.w8(32'h38848e14),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7720ae),
	.w1(32'hbb21f1dd),
	.w2(32'h3b9796f3),
	.w3(32'hbbdcefc4),
	.w4(32'hbb1f287b),
	.w5(32'hbd21f882),
	.w6(32'h3b79130f),
	.w7(32'h3c7b7b69),
	.w8(32'hbca34f36),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3e0208),
	.w1(32'hbb3fa1af),
	.w2(32'h3c1d9b7f),
	.w3(32'hbb185287),
	.w4(32'hbc6df761),
	.w5(32'hbb803bb2),
	.w6(32'h3bfbac9e),
	.w7(32'hbc746ce8),
	.w8(32'h3c1651ca),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b5015),
	.w1(32'hbd8620b4),
	.w2(32'h3b10468e),
	.w3(32'hbb171f73),
	.w4(32'hbab81cc7),
	.w5(32'h3c71ae8f),
	.w6(32'hbb45860a),
	.w7(32'hbb27efa2),
	.w8(32'hbb27edc3),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf370ff),
	.w1(32'h3b36e484),
	.w2(32'hbb373230),
	.w3(32'h3b33fc72),
	.w4(32'hbab09f2e),
	.w5(32'h3b825453),
	.w6(32'hbaf8c5e8),
	.w7(32'hbb7bb726),
	.w8(32'h39583da0),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbada38be),
	.w1(32'h3be310d1),
	.w2(32'hba94d06e),
	.w3(32'h3a98c33b),
	.w4(32'hbc8cee2e),
	.w5(32'hbb83be0d),
	.w6(32'h3c7a8c59),
	.w7(32'h3b73d87d),
	.w8(32'hbb22fb49),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c177d12),
	.w1(32'h3c69ae22),
	.w2(32'hbc907c65),
	.w3(32'h3c9083c7),
	.w4(32'hbd8deca7),
	.w5(32'hbc8f58c8),
	.w6(32'hba95da23),
	.w7(32'hbb3cca04),
	.w8(32'hba720085),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdf70a4),
	.w1(32'h3c0f0b13),
	.w2(32'hbcd724a1),
	.w3(32'hbc7d5e8d),
	.w4(32'h3cd08158),
	.w5(32'h394bdb35),
	.w6(32'hbcafc69e),
	.w7(32'hbb0c9edf),
	.w8(32'h3bb533ad),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4a06cf),
	.w1(32'hbad9b4e8),
	.w2(32'h3bbde700),
	.w3(32'h3a1094b6),
	.w4(32'hba0873aa),
	.w5(32'h3b65c14e),
	.w6(32'hbcdeee7c),
	.w7(32'h3bf1c6cb),
	.w8(32'hbca8415b),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adb30aa),
	.w1(32'h3b5e7168),
	.w2(32'h3b765397),
	.w3(32'h3ae52f8d),
	.w4(32'h3c84f9b6),
	.w5(32'hba292155),
	.w6(32'h3c52579b),
	.w7(32'h3b4afaf4),
	.w8(32'hba5afb7b),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba87ff28),
	.w1(32'h3b9b7221),
	.w2(32'h3c4a8377),
	.w3(32'hba19029e),
	.w4(32'hbb14fef6),
	.w5(32'h3c5f1c6d),
	.w6(32'h3a987a2a),
	.w7(32'hbafcdec5),
	.w8(32'h3997e565),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb001534),
	.w1(32'hbb847e76),
	.w2(32'h3b17e01a),
	.w3(32'hbc5b3403),
	.w4(32'hbc9cead9),
	.w5(32'h3b094a07),
	.w6(32'hbba961fb),
	.w7(32'h3bfbd618),
	.w8(32'h3be0ca8b),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0805b8),
	.w1(32'h3bba4e6a),
	.w2(32'hbc86f371),
	.w3(32'hbc505ba6),
	.w4(32'h3c17976c),
	.w5(32'h3ba7270f),
	.w6(32'hbb8143ab),
	.w7(32'h3b955fcf),
	.w8(32'h3c118d0d),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc49fb7e),
	.w1(32'hbc684d1b),
	.w2(32'hbc466cca),
	.w3(32'h3b89b146),
	.w4(32'hbc269262),
	.w5(32'h3c1f16a2),
	.w6(32'hbab2fb4a),
	.w7(32'h3a477e8b),
	.w8(32'hbb98db91),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1f173c),
	.w1(32'h3d44e3b8),
	.w2(32'hbb927230),
	.w3(32'h3b03c9ea),
	.w4(32'h393304f7),
	.w5(32'hbb9954c0),
	.w6(32'h38b52719),
	.w7(32'h3bd08393),
	.w8(32'h3b88ba90),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3c7323),
	.w1(32'hbb970efc),
	.w2(32'h3b9deef1),
	.w3(32'hbb247da4),
	.w4(32'h3c97a6dd),
	.w5(32'hbda9817f),
	.w6(32'h3b26f4a8),
	.w7(32'h3c5fcaba),
	.w8(32'h3b2f776d),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7ce89b),
	.w1(32'hba3d7b2d),
	.w2(32'hbc214d60),
	.w3(32'h3c0f40dd),
	.w4(32'h3bf05cb7),
	.w5(32'hbb475fd4),
	.w6(32'hbc4b2244),
	.w7(32'h3bff697f),
	.w8(32'hba5b1949),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd420aa),
	.w1(32'hbbfd351b),
	.w2(32'hbbedac3a),
	.w3(32'hbb8ebe2a),
	.w4(32'hbd306e48),
	.w5(32'hbbf23ca6),
	.w6(32'h3c911351),
	.w7(32'h3c203448),
	.w8(32'h3ca99857),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb50eb0),
	.w1(32'hbbcc21f1),
	.w2(32'hbb222f9e),
	.w3(32'hbc01d94f),
	.w4(32'h3c039fa4),
	.w5(32'hbb70fcc0),
	.w6(32'hb902ba8f),
	.w7(32'h3bb4288e),
	.w8(32'h3acc845b),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b95ced0),
	.w1(32'hbb588583),
	.w2(32'hbccaf0ef),
	.w3(32'h3c135d9f),
	.w4(32'h3b2f8ba3),
	.w5(32'h3c19345c),
	.w6(32'hbbab7d42),
	.w7(32'hbc057e45),
	.w8(32'h3a2af6b9),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbfd824),
	.w1(32'h3bed094e),
	.w2(32'h3b89a94f),
	.w3(32'h3aca2456),
	.w4(32'hbb15f291),
	.w5(32'h396980e8),
	.w6(32'hbbbde104),
	.w7(32'hbbb12a04),
	.w8(32'h3bbedba3),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc80820f),
	.w1(32'hbadf07d6),
	.w2(32'hbb8a6850),
	.w3(32'h3d0ed613),
	.w4(32'hbc34a6de),
	.w5(32'hbbd8c1db),
	.w6(32'h3c019dce),
	.w7(32'hbb23e084),
	.w8(32'hbbd1f531),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb44e67c),
	.w1(32'h3b66f26e),
	.w2(32'h3b0b5953),
	.w3(32'hbc662a14),
	.w4(32'hbc574574),
	.w5(32'h3b0d1604),
	.w6(32'hbb1d6ecf),
	.w7(32'h3b912c9f),
	.w8(32'h3cb24658),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bce4132),
	.w1(32'hbd820ecf),
	.w2(32'h3a8da88b),
	.w3(32'hbba75e3b),
	.w4(32'hbbe15c79),
	.w5(32'hbc3878bc),
	.w6(32'h3c0f22ab),
	.w7(32'h3ba6631d),
	.w8(32'hbc91ef30),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c41763c),
	.w1(32'hba5b9311),
	.w2(32'h3be5efaf),
	.w3(32'h3bcd1198),
	.w4(32'hbc5e0a9d),
	.w5(32'hbd010528),
	.w6(32'h3b7cf583),
	.w7(32'h3a1715de),
	.w8(32'hb98b9c0c),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba07615),
	.w1(32'h3b8d86d2),
	.w2(32'hbbfebeba),
	.w3(32'h3aed881e),
	.w4(32'h3b64183d),
	.w5(32'h3c7fc8b0),
	.w6(32'hbc190c34),
	.w7(32'h3a38f44a),
	.w8(32'hbc6c4ba7),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7bda4d),
	.w1(32'hbc7214b5),
	.w2(32'h3be1d468),
	.w3(32'h3bdfd26f),
	.w4(32'hbbe8dd5b),
	.w5(32'h3b9a592b),
	.w6(32'hbac58bb9),
	.w7(32'hba8a7b1c),
	.w8(32'hbc215201),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb09de99),
	.w1(32'h3a32bb84),
	.w2(32'h3caa172c),
	.w3(32'h3c4e560c),
	.w4(32'hba6cdc04),
	.w5(32'hba8a743d),
	.w6(32'h3c24c13a),
	.w7(32'hbb99b9f0),
	.w8(32'h3c32de5c),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93edc4f),
	.w1(32'hbafa2784),
	.w2(32'hbb74881b),
	.w3(32'hbc1d6c67),
	.w4(32'h3beae47c),
	.w5(32'hbac168c5),
	.w6(32'hbb5e6a88),
	.w7(32'h3c0ab470),
	.w8(32'hbbaf93ca),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0f4c2c),
	.w1(32'h3b4259c4),
	.w2(32'hbbae4799),
	.w3(32'hbd171835),
	.w4(32'hbad5020f),
	.w5(32'h3b4c25ed),
	.w6(32'h3c17d1ca),
	.w7(32'hbc0e6c8d),
	.w8(32'hbc162619),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc869521),
	.w1(32'hbc3f4ee1),
	.w2(32'h3b05c85d),
	.w3(32'h3d2e5e1e),
	.w4(32'h3c80ca81),
	.w5(32'h3a3c5b73),
	.w6(32'h3c9b10ea),
	.w7(32'h3985bc0a),
	.w8(32'hbc08b945),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc621093),
	.w1(32'hbb171174),
	.w2(32'hba939d7c),
	.w3(32'h3bf2751d),
	.w4(32'hbc160957),
	.w5(32'hbbf9513f),
	.w6(32'h3bdaf382),
	.w7(32'hb88f1179),
	.w8(32'hbbaff250),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9132ad5),
	.w1(32'h3abbdc12),
	.w2(32'h3c5de9cd),
	.w3(32'hba7dcc43),
	.w4(32'hbc918f30),
	.w5(32'h3c80c4e5),
	.w6(32'h3b0e0849),
	.w7(32'hbc19c964),
	.w8(32'h3c5ce4a7),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb312c35),
	.w1(32'hbc411e54),
	.w2(32'h3c613026),
	.w3(32'h3b82c4cc),
	.w4(32'hbc029baf),
	.w5(32'h3b9297f1),
	.w6(32'hbb984d14),
	.w7(32'hbb360474),
	.w8(32'hbb98cb43),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc0bc9a),
	.w1(32'hb94ec25b),
	.w2(32'h3b50e424),
	.w3(32'h3b98b320),
	.w4(32'h3bee69de),
	.w5(32'hbb302400),
	.w6(32'h3c306d8d),
	.w7(32'h39ee4853),
	.w8(32'h3ba913ee),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7e7d43),
	.w1(32'h3b4685ad),
	.w2(32'hbbbd3624),
	.w3(32'h3bf857c4),
	.w4(32'h3bc40e4b),
	.w5(32'h3c0a5a1d),
	.w6(32'h3b00be6f),
	.w7(32'h3b032e7f),
	.w8(32'h3cd4fe08),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b88c40d),
	.w1(32'hbc4fc785),
	.w2(32'hbbf44162),
	.w3(32'h3b329ce1),
	.w4(32'hbbc910a3),
	.w5(32'h3cc3c43c),
	.w6(32'hbc18f2aa),
	.w7(32'hbc8cb6e9),
	.w8(32'hbc6b99ae),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc86e974),
	.w1(32'hbc8ee38c),
	.w2(32'h3cc40929),
	.w3(32'h3c0cafe5),
	.w4(32'hbc83213a),
	.w5(32'hba518567),
	.w6(32'h3d060f60),
	.w7(32'h3c92fac6),
	.w8(32'h3c612904),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc00939),
	.w1(32'h3c0a4822),
	.w2(32'hb9ba64f8),
	.w3(32'hbc61fd0d),
	.w4(32'hbbadc719),
	.w5(32'hbab567c8),
	.w6(32'h3c1e1e2c),
	.w7(32'h3d3bcd83),
	.w8(32'h3c845c94),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aadf6f8),
	.w1(32'h3c21ddef),
	.w2(32'h3ccccbfd),
	.w3(32'hbb0e28ba),
	.w4(32'h3be25a71),
	.w5(32'hbcbd3c60),
	.w6(32'hbc0eabaf),
	.w7(32'hbbd50d10),
	.w8(32'h3c3b225a),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcbff83),
	.w1(32'hbd237558),
	.w2(32'h3b2ac1e4),
	.w3(32'h3bf4e6f2),
	.w4(32'h3cc0ccca),
	.w5(32'h3b8be6ce),
	.w6(32'h3cc87def),
	.w7(32'hbc37fd75),
	.w8(32'h384aab68),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3badc5bb),
	.w1(32'h3a9b8190),
	.w2(32'hbbd320a1),
	.w3(32'hbbdb84d1),
	.w4(32'hbbf83927),
	.w5(32'h3a806f73),
	.w6(32'h3a900e3e),
	.w7(32'hbc10b1e8),
	.w8(32'h3bbe70d3),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5f2807),
	.w1(32'hbbc2f125),
	.w2(32'h3c04d329),
	.w3(32'h3b1d77c6),
	.w4(32'hbc1b4cc9),
	.w5(32'hbb4b59e3),
	.w6(32'h3bc34df4),
	.w7(32'hbbd52415),
	.w8(32'hba8e17ed),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b83d7f4),
	.w1(32'hbb150041),
	.w2(32'hbc5120b0),
	.w3(32'hba9d215d),
	.w4(32'hbbd69669),
	.w5(32'hb9a26303),
	.w6(32'h3bddab63),
	.w7(32'h3bbe2e16),
	.w8(32'h3c0fd95f),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc510ec8),
	.w1(32'hba484aad),
	.w2(32'h3af0a68b),
	.w3(32'hbbb96ad1),
	.w4(32'hbc3dd726),
	.w5(32'h3b553e04),
	.w6(32'h3a0d3f08),
	.w7(32'hbc36e742),
	.w8(32'h3c09a1a8),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf5c2b4),
	.w1(32'hba4085b2),
	.w2(32'hbc544c48),
	.w3(32'h3bad265a),
	.w4(32'hbc23b811),
	.w5(32'hbae56e39),
	.w6(32'hbb892131),
	.w7(32'hbaa24411),
	.w8(32'h3c5f2e84),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8ab267),
	.w1(32'h3bc2b2f2),
	.w2(32'hbb2a7b2e),
	.w3(32'hbc371c87),
	.w4(32'hbb3169d1),
	.w5(32'hbbd42811),
	.w6(32'h3c596512),
	.w7(32'hba9f8766),
	.w8(32'hbc723f82),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a45a2a4),
	.w1(32'h3b330263),
	.w2(32'hbb121ec3),
	.w3(32'h3aca4e23),
	.w4(32'hbc9ffcf4),
	.w5(32'hbb244874),
	.w6(32'hbbbcfd5e),
	.w7(32'hbc2b1def),
	.w8(32'hbc8718db),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e147ca),
	.w1(32'hbb7f049c),
	.w2(32'hbc33baf9),
	.w3(32'hbb881b43),
	.w4(32'h39753eee),
	.w5(32'hbc196be7),
	.w6(32'hbd016589),
	.w7(32'hbb812b11),
	.w8(32'h3c386911),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b891d1b),
	.w1(32'hbb02df03),
	.w2(32'h3c9b1b2e),
	.w3(32'h3b4aa0aa),
	.w4(32'hbc1ae888),
	.w5(32'hbba51670),
	.w6(32'h38498672),
	.w7(32'hbcc08426),
	.w8(32'h3baeb4f8),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb208b27),
	.w1(32'hbc85a289),
	.w2(32'h3baec455),
	.w3(32'hbb9e68bf),
	.w4(32'hbbf1e3d2),
	.w5(32'h3af5b873),
	.w6(32'hbc84f9aa),
	.w7(32'hbb61277b),
	.w8(32'hbbeedce5),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8cb176),
	.w1(32'h37fc65da),
	.w2(32'h3a21a358),
	.w3(32'hbbe27dea),
	.w4(32'hbc0f6cc4),
	.w5(32'hbb73b425),
	.w6(32'h3c5c67b4),
	.w7(32'h3d0c2e60),
	.w8(32'hbb8ca042),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfa6645),
	.w1(32'hbc70ffec),
	.w2(32'hbaec0807),
	.w3(32'hbb02d243),
	.w4(32'h3c6e02f4),
	.w5(32'hbaae84f2),
	.w6(32'hbbe57ee4),
	.w7(32'h3c96c1f4),
	.w8(32'hbc0b0911),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c91550b),
	.w1(32'hbbbd3f1e),
	.w2(32'hbbde73c3),
	.w3(32'hbbd9efa9),
	.w4(32'h3bb240b2),
	.w5(32'h3b59bcad),
	.w6(32'h3c2a54d7),
	.w7(32'hbca41880),
	.w8(32'hbc5c4d79),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3c5e04),
	.w1(32'hbbf94fd9),
	.w2(32'h3b9e6c9a),
	.w3(32'hbae16625),
	.w4(32'hbc2d7922),
	.w5(32'h3bed1f74),
	.w6(32'h3c1db196),
	.w7(32'h392d637a),
	.w8(32'hbb3dd8c8),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c270d90),
	.w1(32'hba916b55),
	.w2(32'h3b8a600a),
	.w3(32'hba63423c),
	.w4(32'hbbc39eb6),
	.w5(32'h3a413f46),
	.w6(32'h39c7cee3),
	.w7(32'hbc0af2c1),
	.w8(32'hbbb87712),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc62b53),
	.w1(32'h3b80fa3a),
	.w2(32'hbae61127),
	.w3(32'h3c14b851),
	.w4(32'h3a689a32),
	.w5(32'h3b93b69d),
	.w6(32'hbb0f9ee3),
	.w7(32'hbbecdad2),
	.w8(32'h3bcc82ed),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5e10a0),
	.w1(32'hbbf1dab6),
	.w2(32'h3c56b40e),
	.w3(32'hbba97839),
	.w4(32'h3b8e8ac3),
	.w5(32'h3b2b8a4f),
	.w6(32'h3b378bcf),
	.w7(32'hbcb65eb7),
	.w8(32'hbba8e964),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcc469dc),
	.w1(32'hbbca932a),
	.w2(32'h3be4eb2b),
	.w3(32'h3b15078e),
	.w4(32'h39c21468),
	.w5(32'h3bfbf5e4),
	.w6(32'hb8f7fbc7),
	.w7(32'h3c83115f),
	.w8(32'h3c5b1ed1),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1ff35d),
	.w1(32'hbc4b97f1),
	.w2(32'h3c117f1d),
	.w3(32'hbbf055f0),
	.w4(32'hbc3b1a17),
	.w5(32'h3b74a807),
	.w6(32'h3b8c8b41),
	.w7(32'h3c436a5d),
	.w8(32'h3be68a1b),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc164b86),
	.w1(32'hbc019c34),
	.w2(32'h3cb8fe9a),
	.w3(32'h3aa4071f),
	.w4(32'hb8e2b01e),
	.w5(32'hba305a36),
	.w6(32'hba9cee30),
	.w7(32'hbbe45ce4),
	.w8(32'hb84cf3cc),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5db894),
	.w1(32'hbc4d525c),
	.w2(32'hbc173b13),
	.w3(32'h3b989297),
	.w4(32'hbbf5a8cc),
	.w5(32'hbc91fddb),
	.w6(32'h3c04b848),
	.w7(32'hbb190080),
	.w8(32'h3be81f4e),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5a9c1f),
	.w1(32'hbb128353),
	.w2(32'h3ae981e9),
	.w3(32'hba458882),
	.w4(32'h3cb762be),
	.w5(32'hbb89747b),
	.w6(32'hbad70832),
	.w7(32'hbc368a68),
	.w8(32'h3c2d1a10),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad81d2d),
	.w1(32'hbbdd2b53),
	.w2(32'hbc91ef35),
	.w3(32'hbae9645c),
	.w4(32'hbbff8547),
	.w5(32'h3b4b358b),
	.w6(32'h3c1a402e),
	.w7(32'h3ac60fdb),
	.w8(32'h3b836b06),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba16cad),
	.w1(32'h3cc902cc),
	.w2(32'hbb77ad85),
	.w3(32'hbb23f352),
	.w4(32'hbc0b7bc8),
	.w5(32'hbb605a6d),
	.w6(32'hba284f37),
	.w7(32'hbacf314e),
	.w8(32'hbc84deb8),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc70f84e),
	.w1(32'h3aea0388),
	.w2(32'h3c658892),
	.w3(32'hbb1aeb71),
	.w4(32'h3bbe6c7d),
	.w5(32'hbb6fdf2f),
	.w6(32'hbc271b8f),
	.w7(32'h3bf88cc3),
	.w8(32'hbc8168d1),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a81cbf7),
	.w1(32'hbbbd2e55),
	.w2(32'hbb7e3b5e),
	.w3(32'h388971aa),
	.w4(32'hbc3d7608),
	.w5(32'h3c7ed547),
	.w6(32'hbad0a5fb),
	.w7(32'h3ad08c61),
	.w8(32'hb9e29116),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cac04d1),
	.w1(32'h3b897a8d),
	.w2(32'hbbae33ad),
	.w3(32'hbab2af69),
	.w4(32'hbc061261),
	.w5(32'hbb89aa33),
	.w6(32'h3c0e7279),
	.w7(32'h3bb37996),
	.w8(32'hba85cc0b),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5e09c1),
	.w1(32'hbc4d6f5a),
	.w2(32'hbb27bfce),
	.w3(32'h3a12e4ce),
	.w4(32'hbc289f5d),
	.w5(32'hbd640e2b),
	.w6(32'hbd040598),
	.w7(32'h3b65cdd7),
	.w8(32'h3a85361d),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5e1b58),
	.w1(32'hbce392b7),
	.w2(32'hbb14fc44),
	.w3(32'hbc319b73),
	.w4(32'h3b58791c),
	.w5(32'hbcaa56ee),
	.w6(32'h3cbb6ee7),
	.w7(32'hbbc43d32),
	.w8(32'h3c9df464),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc589a4),
	.w1(32'h3c4fd2b1),
	.w2(32'h3b82e240),
	.w3(32'h3bfe38a2),
	.w4(32'h3c4feaee),
	.w5(32'h3bb2c82a),
	.w6(32'hbc07589b),
	.w7(32'hbb4bb3ab),
	.w8(32'hbb982d1b),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc702a83),
	.w1(32'hbafa725b),
	.w2(32'h3c25efa4),
	.w3(32'h3badf5f4),
	.w4(32'h3c0290ba),
	.w5(32'h3b852f62),
	.w6(32'hbb7c8e30),
	.w7(32'h3c054210),
	.w8(32'hbb15c889),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc7a3d6),
	.w1(32'hba5e0bc3),
	.w2(32'hbcbffaff),
	.w3(32'hbc4a8c14),
	.w4(32'hbbb571e5),
	.w5(32'hbc26c0ab),
	.w6(32'hbb115cbb),
	.w7(32'hbc2623d5),
	.w8(32'h3d1cdb47),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb318ddf),
	.w1(32'h3c066889),
	.w2(32'h3c1758ad),
	.w3(32'h3aa72f08),
	.w4(32'hbc13a3d1),
	.w5(32'hbb842a7d),
	.w6(32'hbbdabfbd),
	.w7(32'hbb253cf8),
	.w8(32'h3b8841fd),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a821a01),
	.w1(32'h3c6b9d1c),
	.w2(32'h3c2ee69f),
	.w3(32'hbcba3345),
	.w4(32'hbbf0fbe4),
	.w5(32'hbc9d6075),
	.w6(32'h3bd71631),
	.w7(32'h3ac04fec),
	.w8(32'h3c153460),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1beca7),
	.w1(32'hbc0e1a02),
	.w2(32'h3bcf34d6),
	.w3(32'h3b313f75),
	.w4(32'h3a9fb3d6),
	.w5(32'hbc2e6a72),
	.w6(32'hb8f3b654),
	.w7(32'h3b51b5f9),
	.w8(32'hbc0d6762),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcafa709),
	.w1(32'h3c0c0e47),
	.w2(32'h3c83cb82),
	.w3(32'h3b8ec23f),
	.w4(32'h3b4cfb5f),
	.w5(32'h3bbb6558),
	.w6(32'hbc2a0c63),
	.w7(32'hbcc55fd7),
	.w8(32'h3b9ba019),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3b5c02),
	.w1(32'hbbf09eb5),
	.w2(32'hbb0ce471),
	.w3(32'hbc2f0aa0),
	.w4(32'h3b054ebe),
	.w5(32'h3ae1fcb0),
	.w6(32'h3c61289e),
	.w7(32'h3b596ddb),
	.w8(32'hbc2a386d),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4742ef),
	.w1(32'h3b20e808),
	.w2(32'hbc2dcbdf),
	.w3(32'hbc4fa40d),
	.w4(32'hbbbf813f),
	.w5(32'hbc7d2196),
	.w6(32'hbc492ebd),
	.w7(32'h3c474417),
	.w8(32'h3ca85161),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1276fd),
	.w1(32'hbbfdfed7),
	.w2(32'h3be5f4ad),
	.w3(32'h3afd3ff6),
	.w4(32'hb99e8f4c),
	.w5(32'hbce72c5d),
	.w6(32'h3b7b88f2),
	.w7(32'hbbde3429),
	.w8(32'h3b79732d),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb189356),
	.w1(32'h3c78e66c),
	.w2(32'hbbaf376b),
	.w3(32'h3bcc7105),
	.w4(32'h3c397a73),
	.w5(32'h39f7668c),
	.w6(32'hbc3b9e93),
	.w7(32'hbc30120c),
	.w8(32'hbb1d3543),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb84878),
	.w1(32'hbb9c9aee),
	.w2(32'hbd138062),
	.w3(32'hbbc4e4e2),
	.w4(32'h3bb6f959),
	.w5(32'h3ba2facb),
	.w6(32'hbbf0a9c3),
	.w7(32'h3c11dc28),
	.w8(32'hbbfab33a),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab8ea53),
	.w1(32'h3c3ce27d),
	.w2(32'h3b89dda8),
	.w3(32'hb9a9cace),
	.w4(32'hbbd92762),
	.w5(32'hbbca37cb),
	.w6(32'h3ca9d00b),
	.w7(32'h3cb6babc),
	.w8(32'h3c2732c9),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8ff6af),
	.w1(32'hbc0c9d6c),
	.w2(32'hbbf59d23),
	.w3(32'hbadbc92a),
	.w4(32'hbc5cf1dd),
	.w5(32'hbb772891),
	.w6(32'hbab2bd9d),
	.w7(32'hbba35884),
	.w8(32'hbc6a457e),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc57a85f),
	.w1(32'h3c052a97),
	.w2(32'h39fdcc5f),
	.w3(32'h39457bff),
	.w4(32'hbabc1eac),
	.w5(32'hbddb4797),
	.w6(32'hbc122746),
	.w7(32'hbc1386f8),
	.w8(32'h3c00f7e5),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8b0a6d),
	.w1(32'hbbd434f4),
	.w2(32'hbac5b007),
	.w3(32'hbb937919),
	.w4(32'hbc8077b0),
	.w5(32'h39dd12ca),
	.w6(32'h3c79843e),
	.w7(32'h3b11b417),
	.w8(32'hbb68edbe),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcaad5fe),
	.w1(32'h3c1f6622),
	.w2(32'hbbc78d56),
	.w3(32'hbbaf519f),
	.w4(32'hbc0e1eaa),
	.w5(32'h3c11dabf),
	.w6(32'hbc0f0528),
	.w7(32'hbba25cb5),
	.w8(32'hbcff2a0a),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4a4f38),
	.w1(32'hbbf17441),
	.w2(32'hbc26dcae),
	.w3(32'h3c967853),
	.w4(32'h39b6e3ec),
	.w5(32'h3ad672b1),
	.w6(32'h3b0d2473),
	.w7(32'hbbe9686e),
	.w8(32'h3c7c83ec),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c9cbc13),
	.w1(32'h3ba867f1),
	.w2(32'h3c577925),
	.w3(32'hbb21026d),
	.w4(32'hba17080e),
	.w5(32'h3beda157),
	.w6(32'h3be78c1a),
	.w7(32'h3a688b94),
	.w8(32'h3b26ea3d),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb29b38),
	.w1(32'h3bc50336),
	.w2(32'h3c227cea),
	.w3(32'hbc9ead8b),
	.w4(32'h3c0c6eac),
	.w5(32'hbc4c4bf5),
	.w6(32'hba21945d),
	.w7(32'hb88dca2a),
	.w8(32'hbadccc5d),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc8ed9e),
	.w1(32'h3aa6dfee),
	.w2(32'hbc0ac518),
	.w3(32'hbb3a6955),
	.w4(32'h3a9b64c0),
	.w5(32'hbb6d4f47),
	.w6(32'h3b7b56cd),
	.w7(32'hbc9344dd),
	.w8(32'h3b1e6262),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3c4c60),
	.w1(32'hbabb796c),
	.w2(32'hbccb4e6d),
	.w3(32'h3be9f0ca),
	.w4(32'h3cb2d644),
	.w5(32'hbd18b2ca),
	.w6(32'h3c0d2eb5),
	.w7(32'h3b25e5ce),
	.w8(32'hbaa8f830),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bad6d4b),
	.w1(32'hbac8274c),
	.w2(32'h3c51968c),
	.w3(32'hbcb82036),
	.w4(32'h3c96f87c),
	.w5(32'hbbf5c562),
	.w6(32'hbb9e0dec),
	.w7(32'h3bcc0477),
	.w8(32'h3bffa34c),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b985982),
	.w1(32'h3b9a6ee7),
	.w2(32'h3c3ca1d2),
	.w3(32'h38b1720d),
	.w4(32'hbb540106),
	.w5(32'hbb82e45f),
	.w6(32'hbbdf9616),
	.w7(32'h3c7116ef),
	.w8(32'h3b1f0a02),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bac1f2e),
	.w1(32'h3b85279b),
	.w2(32'hbbef84f0),
	.w3(32'h3c417c71),
	.w4(32'h3c07ebea),
	.w5(32'h3c2b71a5),
	.w6(32'hbc1930fb),
	.w7(32'h3c828c9a),
	.w8(32'h3be66083),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c321637),
	.w1(32'hb8f5bf59),
	.w2(32'h3bcf3d9e),
	.w3(32'h3bada0cc),
	.w4(32'hbcb0de37),
	.w5(32'h3b7cc7ac),
	.w6(32'hbd6ba34c),
	.w7(32'h3ba5c4c6),
	.w8(32'h3c2d5f24),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcfeda2),
	.w1(32'hbb91cc3a),
	.w2(32'hbc29fc3d),
	.w3(32'h3c2e7ca3),
	.w4(32'h3bc80405),
	.w5(32'h3d0242a0),
	.w6(32'h3b5e5b90),
	.w7(32'h3ba47c0d),
	.w8(32'h3ab0de09),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c853d8b),
	.w1(32'hbb9aab4b),
	.w2(32'h398eff48),
	.w3(32'hbcae7f72),
	.w4(32'hbce12a02),
	.w5(32'hbdce0664),
	.w6(32'hbc3382cb),
	.w7(32'h3cfc2219),
	.w8(32'h3ccd5814),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8e7aa6),
	.w1(32'hbcac9f35),
	.w2(32'hbb690720),
	.w3(32'h3ade0ec2),
	.w4(32'h3a9a6a36),
	.w5(32'h3c2ce5b6),
	.w6(32'h3c38a4aa),
	.w7(32'hb9be67c8),
	.w8(32'h3b801c5e),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9fec1f),
	.w1(32'h3b5781b1),
	.w2(32'hbce22663),
	.w3(32'h3b453da9),
	.w4(32'h3b1ca615),
	.w5(32'hbb8b1254),
	.w6(32'hbab5ad37),
	.w7(32'hbbd2715b),
	.w8(32'h3bc503d3),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba96a7c2),
	.w1(32'hbb245d3b),
	.w2(32'h3be5c7fc),
	.w3(32'hbcaef6d2),
	.w4(32'hbc8eee39),
	.w5(32'hbac736a5),
	.w6(32'h3b0a2ee5),
	.w7(32'h3c8c298c),
	.w8(32'h3aaf0db3),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe3f142),
	.w1(32'h3bdedee4),
	.w2(32'h3b008c17),
	.w3(32'hb958d719),
	.w4(32'h3ca6e381),
	.w5(32'hbb1a2dc5),
	.w6(32'hbb72d7ed),
	.w7(32'hbc2edd85),
	.w8(32'hbc0ffb5d),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b960a40),
	.w1(32'hb8b5c85c),
	.w2(32'h3bf6f783),
	.w3(32'h3bfb604e),
	.w4(32'hbb2f0128),
	.w5(32'h3d23faf8),
	.w6(32'h3b3fb576),
	.w7(32'hbd4b6735),
	.w8(32'hbb2f67b3),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0ad2b7),
	.w1(32'hbb848672),
	.w2(32'h3b708c7e),
	.w3(32'hbbaa7d23),
	.w4(32'hbbd90c60),
	.w5(32'h3bd71385),
	.w6(32'hbbbc481c),
	.w7(32'hba1fee49),
	.w8(32'hbbf7f23d),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c73dba7),
	.w1(32'hbc6e4096),
	.w2(32'hbc54541b),
	.w3(32'h39dc122a),
	.w4(32'hbc2679cb),
	.w5(32'h394a1ff0),
	.w6(32'h3bd1947c),
	.w7(32'h3c86d1c1),
	.w8(32'h3895c8cf),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c24dc0e),
	.w1(32'h3a7379dc),
	.w2(32'h3c6df80c),
	.w3(32'h3b7a469a),
	.w4(32'h3bb8205a),
	.w5(32'h3b2b9e4e),
	.w6(32'hbc0c5af0),
	.w7(32'h3aadd3b0),
	.w8(32'hba13eb6e),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7aa62c),
	.w1(32'hba93bdd0),
	.w2(32'hbc047765),
	.w3(32'hba128779),
	.w4(32'hbd0fa78a),
	.w5(32'hbd2de6f6),
	.w6(32'hbb01eabc),
	.w7(32'h3a909558),
	.w8(32'h3c034723),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3969088e),
	.w1(32'hbd9b927b),
	.w2(32'hbb295aa1),
	.w3(32'h3ab3f567),
	.w4(32'hbbb5abdb),
	.w5(32'hbc06b5d8),
	.w6(32'h3c8c057a),
	.w7(32'h3b1821cf),
	.w8(32'h3afdd8ee),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdb9aa6),
	.w1(32'hb9f79d87),
	.w2(32'h3c234692),
	.w3(32'h3c197d76),
	.w4(32'hbc4671b5),
	.w5(32'h3bdc89a5),
	.w6(32'hbc0a2142),
	.w7(32'h3c23cf14),
	.w8(32'hbb29b5a9),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaf962e),
	.w1(32'hbba93784),
	.w2(32'hbbef0c8b),
	.w3(32'hbbedf27c),
	.w4(32'h3bf24652),
	.w5(32'hba853e6f),
	.w6(32'h3c3b8247),
	.w7(32'h3b6e6e92),
	.w8(32'h3bf71244),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab04ede),
	.w1(32'h3a100ed7),
	.w2(32'hbab5b88e),
	.w3(32'hbe1c92d6),
	.w4(32'h3c1745ff),
	.w5(32'hbc383ccb),
	.w6(32'h3aa1f110),
	.w7(32'hbb40680f),
	.w8(32'hbbc9c7cf),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2e3586),
	.w1(32'h3c8ab12c),
	.w2(32'h3ccbe530),
	.w3(32'hbc5e0da1),
	.w4(32'hbc6465fb),
	.w5(32'h3c33859d),
	.w6(32'hbc493fe8),
	.w7(32'h39a0700d),
	.w8(32'hbc116b60),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc13dd8),
	.w1(32'hbb299aa7),
	.w2(32'h3c3e5e97),
	.w3(32'hbb828c30),
	.w4(32'hbc2d7184),
	.w5(32'h3c308c87),
	.w6(32'h3ae81e58),
	.w7(32'hbbf6a4b7),
	.w8(32'hbadb9fe8),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c410b61),
	.w1(32'hbc01b4bf),
	.w2(32'h3b0a00f0),
	.w3(32'h3b1e77bb),
	.w4(32'hbb88187f),
	.w5(32'hbb2a6979),
	.w6(32'h3c85628c),
	.w7(32'hbb763866),
	.w8(32'h3b225835),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb75b875),
	.w1(32'hbc1f45bc),
	.w2(32'h3b4541b7),
	.w3(32'hbb2c8645),
	.w4(32'h3c818989),
	.w5(32'h3c5283be),
	.w6(32'hbab9997c),
	.w7(32'h3bb68911),
	.w8(32'h3b1f91bd),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b26ed52),
	.w1(32'h3c8d49d6),
	.w2(32'hbb9f5f40),
	.w3(32'hbb21dafa),
	.w4(32'hbb08b0f7),
	.w5(32'h3bd85029),
	.w6(32'h3b6b692e),
	.w7(32'h3ba560ad),
	.w8(32'hbb1de811),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae593ef),
	.w1(32'hbd22b31e),
	.w2(32'h3c4e54e8),
	.w3(32'h3b416a76),
	.w4(32'h3c00b9ea),
	.w5(32'h3ae1c54a),
	.w6(32'h3ba6a329),
	.w7(32'hbc23819c),
	.w8(32'h3b979e1a),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a46b374),
	.w1(32'h3afa7e63),
	.w2(32'h3ba14598),
	.w3(32'hbcc93e77),
	.w4(32'hbc6cbb6b),
	.w5(32'hb9102896),
	.w6(32'hbbaca39e),
	.w7(32'hbd130fd1),
	.w8(32'h3add3010),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2df058),
	.w1(32'hbca4d0da),
	.w2(32'h3c205898),
	.w3(32'h3c2d5254),
	.w4(32'h39d8d0a7),
	.w5(32'hbabe8b25),
	.w6(32'hbb79346d),
	.w7(32'hbbc3b093),
	.w8(32'hbae8325a),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb85af49),
	.w1(32'h3c26b012),
	.w2(32'hbc416932),
	.w3(32'hbc1649ee),
	.w4(32'h3b304b9d),
	.w5(32'hbbe83ac6),
	.w6(32'hbb8b05a1),
	.w7(32'hbb0ae6b9),
	.w8(32'h3a1ab033),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb785206c),
	.w1(32'h3bee27b9),
	.w2(32'hbc751d16),
	.w3(32'h3a8f6559),
	.w4(32'hbc547e07),
	.w5(32'h3b97c696),
	.w6(32'h3b174daa),
	.w7(32'h39e4dc98),
	.w8(32'hbc3972a4),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b830642),
	.w1(32'hb9162bad),
	.w2(32'hbc3be8e2),
	.w3(32'h3bd3e266),
	.w4(32'hbc009e0a),
	.w5(32'h3b5312f3),
	.w6(32'hbc437a32),
	.w7(32'hbb89bb48),
	.w8(32'hbc301e7a),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb060ad),
	.w1(32'h3b733bb8),
	.w2(32'h3b150cf3),
	.w3(32'hbc31cc6c),
	.w4(32'hbb450b66),
	.w5(32'h3c70ec36),
	.w6(32'hbb961862),
	.w7(32'hbc500dc0),
	.w8(32'h3b655963),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc9a9618),
	.w1(32'h3ba4ae17),
	.w2(32'h3c017e86),
	.w3(32'hbc004aed),
	.w4(32'hba90dbd4),
	.w5(32'h39344994),
	.w6(32'h3c37465d),
	.w7(32'hba4a4e33),
	.w8(32'hbbdfcce2),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af7104a),
	.w1(32'h3965fd5d),
	.w2(32'hbb51cca3),
	.w3(32'hbb711b04),
	.w4(32'h3c116269),
	.w5(32'hba187677),
	.w6(32'h3bb79b77),
	.w7(32'h3ba1faa5),
	.w8(32'h3c0376f5),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f494a2),
	.w1(32'h3c0c5e6d),
	.w2(32'hbb0db37b),
	.w3(32'hbb96201a),
	.w4(32'h3b594d6f),
	.w5(32'h3bc52870),
	.w6(32'hbc1d8976),
	.w7(32'hbb6265ce),
	.w8(32'h3b2bc9f9),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6495c5),
	.w1(32'h386ed7d3),
	.w2(32'hbbd745ee),
	.w3(32'h3be13417),
	.w4(32'h3c8b8be4),
	.w5(32'h3b77f3c8),
	.w6(32'h397cb539),
	.w7(32'hbab62f4a),
	.w8(32'hba35e837),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bce76c6),
	.w1(32'h3b85203e),
	.w2(32'hbaceee8e),
	.w3(32'h397f6e92),
	.w4(32'hbb67d21b),
	.w5(32'h3c1a0201),
	.w6(32'hbbd1f4cc),
	.w7(32'hbaa806a2),
	.w8(32'h3a8ab734),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0b9da8),
	.w1(32'hbb5ca3f2),
	.w2(32'hbaf36f87),
	.w3(32'hbcd8c3df),
	.w4(32'h3a271d95),
	.w5(32'hba2edb79),
	.w6(32'h3c1b844a),
	.w7(32'hbc4cfe38),
	.w8(32'hbab8c3fe),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8c6cd4),
	.w1(32'h3c2603e7),
	.w2(32'hbcab3c9f),
	.w3(32'hbb569d84),
	.w4(32'h3c88e3ba),
	.w5(32'hbd7b7284),
	.w6(32'h3b79c2cc),
	.w7(32'h3c62bc7b),
	.w8(32'hbad68039),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a5e721),
	.w1(32'h3b1ce2bb),
	.w2(32'h3a5c8c3d),
	.w3(32'h3c498dc9),
	.w4(32'hbc54e764),
	.w5(32'hbbe8d6d9),
	.w6(32'h3b50c96e),
	.w7(32'h3c6314da),
	.w8(32'h3c15af56),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6f2c1f),
	.w1(32'h3c1dc62d),
	.w2(32'h3ce2a5c7),
	.w3(32'h3bd2dba4),
	.w4(32'h3b361832),
	.w5(32'h3bbef849),
	.w6(32'h3c948b48),
	.w7(32'h3b966e78),
	.w8(32'h3c4d1961),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8fced1),
	.w1(32'h3b8217d5),
	.w2(32'h3b377434),
	.w3(32'hbca5d524),
	.w4(32'h39729aa5),
	.w5(32'h3b847d78),
	.w6(32'h3b791254),
	.w7(32'h3bf2ba4a),
	.w8(32'h3c9cce52),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cc90a5),
	.w1(32'hbba0ef72),
	.w2(32'h3af36666),
	.w3(32'hbc6562b9),
	.w4(32'hbd6bb619),
	.w5(32'h3b2cd715),
	.w6(32'hbc4f0830),
	.w7(32'h3bfadc70),
	.w8(32'h3afd3382),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9c89b5),
	.w1(32'h3a057e22),
	.w2(32'hb9951468),
	.w3(32'h3ab37011),
	.w4(32'hbab06842),
	.w5(32'hbb9433d0),
	.w6(32'h3bc3252c),
	.w7(32'h3bc424cf),
	.w8(32'hbcaf9fac),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c684945),
	.w1(32'hba230cdf),
	.w2(32'h39cc299c),
	.w3(32'hbc8277f6),
	.w4(32'h3bc3110e),
	.w5(32'h3c42b0ec),
	.w6(32'hbcc64be3),
	.w7(32'h3ad959aa),
	.w8(32'h3b5d0360),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb96904d),
	.w1(32'hb9ba02ae),
	.w2(32'hbd10e37c),
	.w3(32'hbb987fa6),
	.w4(32'h3bac3d51),
	.w5(32'hbbb48ff3),
	.w6(32'hbae10f8c),
	.w7(32'hb9d4f9f6),
	.w8(32'h3b1f3e42),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9406f0),
	.w1(32'h3b0d68ae),
	.w2(32'h3a98630b),
	.w3(32'hbd0f5600),
	.w4(32'hbae39d02),
	.w5(32'h39db8ec0),
	.w6(32'hba9aa517),
	.w7(32'hbb15029b),
	.w8(32'h3ab35915),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ee3d8d),
	.w1(32'hbbfff12c),
	.w2(32'hba86a7ef),
	.w3(32'h3c458d12),
	.w4(32'h3bc8628b),
	.w5(32'h3aa92d68),
	.w6(32'h3d0a2ebb),
	.w7(32'h3c3b134a),
	.w8(32'h3bd0ed6d),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2ee4a1),
	.w1(32'h3cab53dc),
	.w2(32'h3bc619db),
	.w3(32'hbb8283fc),
	.w4(32'h3ba4530b),
	.w5(32'hbcaca434),
	.w6(32'hbbc0e5f6),
	.w7(32'h3b83d696),
	.w8(32'hba4defef),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcc3d5a),
	.w1(32'hbaccabc5),
	.w2(32'h3b97fc4c),
	.w3(32'hbb680f1c),
	.w4(32'h3abcd03a),
	.w5(32'h3b552f1d),
	.w6(32'h392c641b),
	.w7(32'hbb7e6c71),
	.w8(32'hbbb244ab),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcf40df),
	.w1(32'h3c115f4f),
	.w2(32'h3bedcc5f),
	.w3(32'hbb213f2d),
	.w4(32'hbc13811b),
	.w5(32'h3c2dc153),
	.w6(32'hb978672e),
	.w7(32'hbaeb022c),
	.w8(32'hbc1b5e1c),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe52e0b),
	.w1(32'h3d524a19),
	.w2(32'h3ad0a536),
	.w3(32'h3adb6d89),
	.w4(32'hbc12abea),
	.w5(32'h3c148b8d),
	.w6(32'hbbb1e4c2),
	.w7(32'hbb94d375),
	.w8(32'h3c35b9ac),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe1e030),
	.w1(32'h3b9baa45),
	.w2(32'h3a049584),
	.w3(32'hbc446ea0),
	.w4(32'h3b445da1),
	.w5(32'hbc2ed3c5),
	.w6(32'h3bbcf886),
	.w7(32'hbc6f756a),
	.w8(32'hbaa85ea2),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc871e93),
	.w1(32'h3bde9ee6),
	.w2(32'h3b5b2889),
	.w3(32'hbc25bd90),
	.w4(32'hbb0cfd85),
	.w5(32'h3aae22f5),
	.w6(32'h3c44fb9b),
	.w7(32'h3bb0a2be),
	.w8(32'h3b38cbbb),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6a35e1),
	.w1(32'h3a5f1e24),
	.w2(32'h3bafca55),
	.w3(32'h3b78dc50),
	.w4(32'hbb3ccce6),
	.w5(32'h3b83990e),
	.w6(32'h3abecb96),
	.w7(32'h3d3e8fa8),
	.w8(32'hbb086d4c),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7b61b7),
	.w1(32'hbc2d79e5),
	.w2(32'h3aa19bec),
	.w3(32'h3bfd8743),
	.w4(32'h3bf6d732),
	.w5(32'h3b239a09),
	.w6(32'hbc7c50f3),
	.w7(32'h3a59f0ba),
	.w8(32'hbb8ed5e7),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0c0ff2),
	.w1(32'h3bdbfde7),
	.w2(32'h3c138875),
	.w3(32'hbc70848c),
	.w4(32'hbce25787),
	.w5(32'hbb7ea4c6),
	.w6(32'h3b2b1946),
	.w7(32'hbca8a9d0),
	.w8(32'h3c96ced5),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9cab21),
	.w1(32'hba290e23),
	.w2(32'h3c7c26e5),
	.w3(32'h3c1e4323),
	.w4(32'hbad6c962),
	.w5(32'hbbbc8642),
	.w6(32'h3baf892b),
	.w7(32'hbbd9656e),
	.w8(32'h3bcce893),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c33d617),
	.w1(32'hbc99923d),
	.w2(32'hbb6502ec),
	.w3(32'hbb1a7a23),
	.w4(32'hb8dab412),
	.w5(32'h3a928002),
	.w6(32'h3bcaa48f),
	.w7(32'h3b19cdf6),
	.w8(32'hbc420cde),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b15fda8),
	.w1(32'hbaa3427d),
	.w2(32'hbbc36239),
	.w3(32'h3b522279),
	.w4(32'hbc53687c),
	.w5(32'hbb3dd9c3),
	.w6(32'hbc7b5c05),
	.w7(32'hbc7e6b5d),
	.w8(32'hbb0ab84c),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdccb0c),
	.w1(32'h3b41e953),
	.w2(32'hbb1399ab),
	.w3(32'h3b648704),
	.w4(32'hbc25b28f),
	.w5(32'hbb8a581a),
	.w6(32'hbc097d49),
	.w7(32'hbbcc11d2),
	.w8(32'h3bbea9f1),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb283da5),
	.w1(32'h3c975641),
	.w2(32'hbc16ab16),
	.w3(32'hbc4da9f3),
	.w4(32'h3b272391),
	.w5(32'hbbd648b9),
	.w6(32'h3a6c27af),
	.w7(32'hbcaa48c5),
	.w8(32'h3bbb0c8c),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1c76a1),
	.w1(32'h3bab418f),
	.w2(32'h3cba5501),
	.w3(32'hbba386c7),
	.w4(32'hbb56e9ad),
	.w5(32'hbb285ee6),
	.w6(32'hbc27617a),
	.w7(32'h3cd1be5d),
	.w8(32'hbc151ff7),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb563d5d),
	.w1(32'hbbe3428c),
	.w2(32'hbc86c4cb),
	.w3(32'hba4641f6),
	.w4(32'h3c82e5c1),
	.w5(32'h3b2ef2f4),
	.w6(32'hbc160943),
	.w7(32'hbca5cb40),
	.w8(32'h3c110e07),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c05a838),
	.w1(32'h3b2ac778),
	.w2(32'hbc19a370),
	.w3(32'hbcc8dc35),
	.w4(32'hbbd01442),
	.w5(32'hbcc8dea4),
	.w6(32'hbada211f),
	.w7(32'h3b2cdb16),
	.w8(32'h3c26ea2a),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcbd13f),
	.w1(32'hbc0d054f),
	.w2(32'hb9df7b2d),
	.w3(32'h3b83c5e2),
	.w4(32'h3aa91f8c),
	.w5(32'h3ba847a5),
	.w6(32'hbbb64037),
	.w7(32'h3d047d5a),
	.w8(32'hbae2df13),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc03b1c0),
	.w1(32'hbc0927b8),
	.w2(32'h3aac3959),
	.w3(32'hb949fe51),
	.w4(32'hbbcf4ea7),
	.w5(32'h3abe2a6c),
	.w6(32'h3c7bbe36),
	.w7(32'h3c1ac73f),
	.w8(32'h3c1c98c5),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d783c22),
	.w1(32'hbc922ddc),
	.w2(32'hbbb68254),
	.w3(32'hbce8efd8),
	.w4(32'h3c420a9f),
	.w5(32'h3c594eb3),
	.w6(32'hbc43e62b),
	.w7(32'hbc33bdca),
	.w8(32'hbc1767ca),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389b0afc),
	.w1(32'hbaa19ec0),
	.w2(32'hbbce7238),
	.w3(32'hbc06a4c8),
	.w4(32'hbc3ba5a7),
	.w5(32'hbb600745),
	.w6(32'hbbd966fd),
	.w7(32'hbb4cd5ef),
	.w8(32'hbc72b1be),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb59aea3),
	.w1(32'h3ba193dd),
	.w2(32'hbc2f23c3),
	.w3(32'hbb87d6f2),
	.w4(32'hba9788c5),
	.w5(32'h3c2766ee),
	.w6(32'h3c31fe92),
	.w7(32'hb92d6f17),
	.w8(32'h3b67b4c8),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2e7aa6),
	.w1(32'h3b07d73d),
	.w2(32'hbd03528a),
	.w3(32'hbb21c9e3),
	.w4(32'h380af976),
	.w5(32'h3b9789fa),
	.w6(32'hbab20b1e),
	.w7(32'h3cc20601),
	.w8(32'h3bdf7741),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6a641c),
	.w1(32'hbbe80c13),
	.w2(32'h399c84f9),
	.w3(32'h399d367d),
	.w4(32'hbc81f478),
	.w5(32'hbb99a2c5),
	.w6(32'hba1977b3),
	.w7(32'hbaceb492),
	.w8(32'h3abd8048),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38175ac9),
	.w1(32'hbc9ae369),
	.w2(32'h3d282eb2),
	.w3(32'hbb902b1d),
	.w4(32'h3cf0383e),
	.w5(32'hbc4a10fd),
	.w6(32'h3c06b2c3),
	.w7(32'hbab12074),
	.w8(32'h3c0716c1),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3452c0),
	.w1(32'h3b199e1d),
	.w2(32'h3cb775e2),
	.w3(32'h3b814891),
	.w4(32'h3ba21dfa),
	.w5(32'hbbe80ab0),
	.w6(32'h3d075f6d),
	.w7(32'hbbb62af5),
	.w8(32'h3b24b590),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2ad019),
	.w1(32'h3b63ea46),
	.w2(32'hbb2faafc),
	.w3(32'hbcc2df8a),
	.w4(32'h3b236c04),
	.w5(32'hbbfbafba),
	.w6(32'hbbacb287),
	.w7(32'hbc791857),
	.w8(32'h3954b0f1),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5c5e25),
	.w1(32'h3bce5408),
	.w2(32'hb8021db2),
	.w3(32'hbb6bc6d9),
	.w4(32'hbb7965d8),
	.w5(32'hbb87eae7),
	.w6(32'h3b779e23),
	.w7(32'h3b25b052),
	.w8(32'hba035ee3),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cfc89b2),
	.w1(32'hbc447e5b),
	.w2(32'hbb7a1caf),
	.w3(32'hbc09c519),
	.w4(32'hbbe0f3e0),
	.w5(32'h3a7fadee),
	.w6(32'hbbdcb857),
	.w7(32'h3b163234),
	.w8(32'h3a6af142),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaf0790),
	.w1(32'h3a675816),
	.w2(32'hba400a05),
	.w3(32'hbb381f66),
	.w4(32'h3c5ebff9),
	.w5(32'h3b05ed22),
	.w6(32'hbbc48d7b),
	.w7(32'hbaeb945a),
	.w8(32'h3c203292),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc20bb4d),
	.w1(32'h3d1454d9),
	.w2(32'h3bc39145),
	.w3(32'h3be5885b),
	.w4(32'h3b956600),
	.w5(32'h3ad2e2a9),
	.w6(32'h3a8f3d3a),
	.w7(32'hbae5c488),
	.w8(32'h3c758505),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba94bac),
	.w1(32'hbc0a37f8),
	.w2(32'hbc667f3b),
	.w3(32'hbbb4231e),
	.w4(32'hbbee5d2c),
	.w5(32'h3c934fbc),
	.w6(32'hbb3caad8),
	.w7(32'hbb20e144),
	.w8(32'hba379420),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a298fe1),
	.w1(32'hbd25b5c9),
	.w2(32'hbbef286e),
	.w3(32'h3bf3a5ec),
	.w4(32'hbbcb280e),
	.w5(32'h3b340bd1),
	.w6(32'h3bb18438),
	.w7(32'h3c11e75a),
	.w8(32'h3c488abb),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdb776e),
	.w1(32'h3ab3e0fc),
	.w2(32'h3c0df72b),
	.w3(32'h3bb9924d),
	.w4(32'hbd09cf3f),
	.w5(32'hbb65e55f),
	.w6(32'h3c5a5301),
	.w7(32'h3bc86d3c),
	.w8(32'hbbf84f46),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3babee13),
	.w1(32'hbc657786),
	.w2(32'hbba664fb),
	.w3(32'hbc11053e),
	.w4(32'hbc195c29),
	.w5(32'h3b9b3dea),
	.w6(32'hbd103f8a),
	.w7(32'h3b855287),
	.w8(32'hba419b39),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbda3d835),
	.w1(32'hbc4dcf43),
	.w2(32'hbb3e625c),
	.w3(32'hbb9481b1),
	.w4(32'h3b1095f3),
	.w5(32'h3b361d0b),
	.w6(32'hbbb8cca7),
	.w7(32'hb90bd850),
	.w8(32'h3b7ce0c2),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aadb048),
	.w1(32'hbba8e786),
	.w2(32'h3bac2750),
	.w3(32'h3a28e898),
	.w4(32'hbb682993),
	.w5(32'h3c063639),
	.w6(32'h3b5a053f),
	.w7(32'h3c9e05ad),
	.w8(32'h3c858a33),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2dca33),
	.w1(32'hbc400264),
	.w2(32'h3a73a76f),
	.w3(32'hbc05451a),
	.w4(32'h3b652c38),
	.w5(32'h3bcf5fbe),
	.w6(32'hba56ce1f),
	.w7(32'h3b1a087a),
	.w8(32'h3ba31142),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7fb3af),
	.w1(32'hbca7f483),
	.w2(32'hba00d205),
	.w3(32'hbc2d3689),
	.w4(32'hb985f6b6),
	.w5(32'h3cada835),
	.w6(32'hbb6dad8c),
	.w7(32'hbba9c5a3),
	.w8(32'h3b1db566),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398cc31a),
	.w1(32'hbce03531),
	.w2(32'h3c2a60da),
	.w3(32'h3cbb7f52),
	.w4(32'hbbb3f5e9),
	.w5(32'h3bd6c0b3),
	.w6(32'h3ab44abe),
	.w7(32'h3c6a147a),
	.w8(32'h3af22454),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb54a7d),
	.w1(32'hba41b43e),
	.w2(32'hbb2079da),
	.w3(32'hbb51ef3b),
	.w4(32'hbc382464),
	.w5(32'h3af31e11),
	.w6(32'hbbc6774c),
	.w7(32'h3b905236),
	.w8(32'h3b08aeba),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb315dd0),
	.w1(32'h386f2dfe),
	.w2(32'h3a23725e),
	.w3(32'hba9de5f3),
	.w4(32'h3bb626b1),
	.w5(32'h3b609525),
	.w6(32'h3bc554b6),
	.w7(32'h3b51f865),
	.w8(32'hb838433a),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a4081),
	.w1(32'hbab5db55),
	.w2(32'hbb6b63d8),
	.w3(32'h3c02b198),
	.w4(32'h3b26cf2c),
	.w5(32'hbc496f85),
	.w6(32'h3c407542),
	.w7(32'h3c3b3bd9),
	.w8(32'h3c4d21b4),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca1ba8d),
	.w1(32'h3bb7242a),
	.w2(32'h39f77f3b),
	.w3(32'h3c2a79d3),
	.w4(32'h3be9fbdc),
	.w5(32'h3a23f88c),
	.w6(32'h3bb56592),
	.w7(32'hbc86add3),
	.w8(32'h3c6ae95f),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6872d4),
	.w1(32'hbba2ef8b),
	.w2(32'h3bff214d),
	.w3(32'hbc92051e),
	.w4(32'h3b9b538b),
	.w5(32'hbb661c06),
	.w6(32'hb92588d0),
	.w7(32'hbb316ad9),
	.w8(32'hbb46f01c),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba21b419),
	.w1(32'hba29151c),
	.w2(32'hbc9a02ff),
	.w3(32'hbb5bf1b3),
	.w4(32'h3b1fc43a),
	.w5(32'h3c505b60),
	.w6(32'h3c4516bf),
	.w7(32'hba9cdcb4),
	.w8(32'hbc1f1494),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8a6722),
	.w1(32'hbc2d3716),
	.w2(32'hbb66fb0b),
	.w3(32'h3a22cd4a),
	.w4(32'hbc437244),
	.w5(32'hbb70a1a2),
	.w6(32'hbade564d),
	.w7(32'h3ade89db),
	.w8(32'hbbb66f2f),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e6d592),
	.w1(32'h3c255039),
	.w2(32'hbd040376),
	.w3(32'h3befa4c0),
	.w4(32'hbc4fdcbd),
	.w5(32'hbb6b00ce),
	.w6(32'hbb49d16a),
	.w7(32'h3c896d70),
	.w8(32'h3bd9a6de),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3ff594),
	.w1(32'hbc3f0185),
	.w2(32'hbc6c5ad5),
	.w3(32'hb93f0d1c),
	.w4(32'hbcb651d5),
	.w5(32'hbc2d4159),
	.w6(32'h3b849051),
	.w7(32'h3b043267),
	.w8(32'h3c83223f),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba153866),
	.w1(32'hbc0da568),
	.w2(32'hbbf6cd27),
	.w3(32'hbcb5a082),
	.w4(32'hbc32fc72),
	.w5(32'hbbf7ce08),
	.w6(32'h3c7b85b2),
	.w7(32'h3d8df75e),
	.w8(32'h3c894211),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9411b8),
	.w1(32'hbc187318),
	.w2(32'hbbf1dc1e),
	.w3(32'h3b95d961),
	.w4(32'hbbaf40af),
	.w5(32'h3ce03b53),
	.w6(32'h3b2f69ee),
	.w7(32'h3c049a54),
	.w8(32'h3be7019c),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb4c213),
	.w1(32'h3bc48cb7),
	.w2(32'h3ba06f8f),
	.w3(32'hbcff1f5b),
	.w4(32'hbb0c00da),
	.w5(32'hbab6aa8d),
	.w6(32'hbb618601),
	.w7(32'hbb342fd0),
	.w8(32'hbc286ca8),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb42b02e),
	.w1(32'h3b378869),
	.w2(32'hbb4c1fb8),
	.w3(32'hba3fd25a),
	.w4(32'h3b22f5c5),
	.w5(32'h3d06c07d),
	.w6(32'hbc2e6c1a),
	.w7(32'hbb911f39),
	.w8(32'h3c83f9ac),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c037b49),
	.w1(32'h3afe0295),
	.w2(32'hbba59d23),
	.w3(32'hbbff7138),
	.w4(32'hbb158bca),
	.w5(32'hbb6a00ff),
	.w6(32'h3b1d118c),
	.w7(32'hbbd96dd7),
	.w8(32'hbb1bd4da),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a53e4fb),
	.w1(32'h386540ce),
	.w2(32'h3c3d6d65),
	.w3(32'hb97fa79e),
	.w4(32'hbb641c3f),
	.w5(32'h3948e0a8),
	.w6(32'h3b80fbd4),
	.w7(32'hbb2b9eeb),
	.w8(32'hbc1dbba9),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca0a95b),
	.w1(32'h3b53dafc),
	.w2(32'h3c199208),
	.w3(32'hbc9371f9),
	.w4(32'hb9755f71),
	.w5(32'h3b2dde23),
	.w6(32'h3c9db2c9),
	.w7(32'hbc1f5b7a),
	.w8(32'h3a71973d),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc07430f),
	.w1(32'hbb7d93da),
	.w2(32'h396fe78e),
	.w3(32'hbb3450b8),
	.w4(32'h3c821d8f),
	.w5(32'h3b6c3bee),
	.w6(32'hbbc34b2f),
	.w7(32'hbb49164d),
	.w8(32'h3aaa1a73),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb1e282),
	.w1(32'hbb8c7451),
	.w2(32'hbc0b9748),
	.w3(32'h3a431a8d),
	.w4(32'hbb8db63a),
	.w5(32'hbd069fdf),
	.w6(32'hbc083080),
	.w7(32'hba04941e),
	.w8(32'h3bb4090a),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3cc734),
	.w1(32'hbc808299),
	.w2(32'hba9a7802),
	.w3(32'h3b35c7eb),
	.w4(32'hb92ecf9b),
	.w5(32'hbbdbb674),
	.w6(32'h3b26c5af),
	.w7(32'h3bf36f3b),
	.w8(32'h3b958153),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b680f),
	.w1(32'h3c8db93b),
	.w2(32'hba2c9365),
	.w3(32'hbb837597),
	.w4(32'hbb08e847),
	.w5(32'hbc0f8c9f),
	.w6(32'h39bb4d50),
	.w7(32'h3c34cae2),
	.w8(32'hbb855b92),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c22b57a),
	.w1(32'hbbd22c23),
	.w2(32'h3c04655e),
	.w3(32'hbc27ad0d),
	.w4(32'hbb429b13),
	.w5(32'h3a92c885),
	.w6(32'hbc9fbc91),
	.w7(32'h3bc32f9d),
	.w8(32'h39801ad9),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4bf842),
	.w1(32'hbc1a735f),
	.w2(32'hbc972f27),
	.w3(32'hbc1d7e97),
	.w4(32'hbc2c55a1),
	.w5(32'hbc7454cd),
	.w6(32'h3bbec015),
	.w7(32'h3b41eb42),
	.w8(32'h3d2e2568),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbafdc6),
	.w1(32'hb9b2c8cb),
	.w2(32'h3b8daca7),
	.w3(32'hbbd0fdf0),
	.w4(32'h3a8b8128),
	.w5(32'h3c51215e),
	.w6(32'hb8b02e25),
	.w7(32'hbb04ab68),
	.w8(32'h3c0374c2),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb78bfe5b),
	.w1(32'h3b37bb44),
	.w2(32'hbb98af0b),
	.w3(32'h3982a6a4),
	.w4(32'h3d118104),
	.w5(32'h3a461282),
	.w6(32'h3a810e39),
	.w7(32'h3b8d868f),
	.w8(32'h3beab175),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab15e9e),
	.w1(32'hbbfcb31b),
	.w2(32'hbcbb6e39),
	.w3(32'hbb2eaffb),
	.w4(32'hbaf15bb6),
	.w5(32'hbb167857),
	.w6(32'h3c4b0683),
	.w7(32'hbb20348a),
	.w8(32'h3ac61885),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd583ed3),
	.w1(32'h3c41d74a),
	.w2(32'h3b51184a),
	.w3(32'h3b8bb3e5),
	.w4(32'hbbd80f21),
	.w5(32'hbc012570),
	.w6(32'h3a27b950),
	.w7(32'hbbb13f6c),
	.w8(32'h3c7f32dd),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc521d96),
	.w1(32'h3b0a3ec0),
	.w2(32'h3c3090dd),
	.w3(32'h3c46f0c0),
	.w4(32'hbc1f6299),
	.w5(32'hbbac786c),
	.w6(32'h3bb2db29),
	.w7(32'h3afec318),
	.w8(32'h3c8dafba),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3ba64b),
	.w1(32'h3c0e84ab),
	.w2(32'hb9d18043),
	.w3(32'hbb6295ac),
	.w4(32'h3bb6f7ed),
	.w5(32'h3cbf502d),
	.w6(32'h3c7575c7),
	.w7(32'hbbf4437d),
	.w8(32'hbb25e61d),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cd4673),
	.w1(32'hbb418076),
	.w2(32'h3c5b66ec),
	.w3(32'hbc28ec5b),
	.w4(32'h3ad4f177),
	.w5(32'h3ae9ad05),
	.w6(32'h3bd8af86),
	.w7(32'hbc1f715a),
	.w8(32'hbc0ae70d),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc960551),
	.w1(32'hbb6d4916),
	.w2(32'h3ad99280),
	.w3(32'h3a479a92),
	.w4(32'h3beeb46a),
	.w5(32'h3bdd3fd0),
	.w6(32'h3a7cf528),
	.w7(32'hb9475b87),
	.w8(32'h3a856b6f),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd3ef38d),
	.w1(32'hbbb876f7),
	.w2(32'hbae93a9d),
	.w3(32'hbaaf0946),
	.w4(32'hbb013f2d),
	.w5(32'h3c7bcd63),
	.w6(32'hbcaf5ba2),
	.w7(32'hbbf97a8b),
	.w8(32'hb899d945),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb95c12f),
	.w1(32'h3c1b1fbe),
	.w2(32'h3b64717f),
	.w3(32'h38bfcef4),
	.w4(32'hbc20818a),
	.w5(32'h3ccf024f),
	.w6(32'h3b2a17c4),
	.w7(32'h3bfbec40),
	.w8(32'hbbab7a0e),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd81237),
	.w1(32'hbce2da03),
	.w2(32'hbc3f70ba),
	.w3(32'hbbbf440e),
	.w4(32'h3c2b3ead),
	.w5(32'hbaa44ce2),
	.w6(32'h3c259133),
	.w7(32'hbc04b7fe),
	.w8(32'hbb512481),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd15602),
	.w1(32'h3b093046),
	.w2(32'h3a6d16f6),
	.w3(32'h3b7a95ee),
	.w4(32'h3afe2684),
	.w5(32'hbb8d6b8e),
	.w6(32'h3b98f83f),
	.w7(32'h3a908638),
	.w8(32'hbbb1ba3e),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2fa664),
	.w1(32'hb9e54da2),
	.w2(32'h39687744),
	.w3(32'hbbf83569),
	.w4(32'h3c681afe),
	.w5(32'h3b79d71b),
	.w6(32'h3adc19aa),
	.w7(32'hbb2c28e3),
	.w8(32'h3bfc1eab),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab714f0),
	.w1(32'hbc43e72d),
	.w2(32'h3b2cf5de),
	.w3(32'h3b5a8585),
	.w4(32'h3aafff26),
	.w5(32'h3c0d5498),
	.w6(32'h3b39560d),
	.w7(32'h3b18594a),
	.w8(32'hbb6c398e),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e05b1),
	.w1(32'h3b9d3c9a),
	.w2(32'h3ab7b9b4),
	.w3(32'h3cf75e8d),
	.w4(32'hbc406b0b),
	.w5(32'hbc6971d3),
	.w6(32'hbc2e7b61),
	.w7(32'h3bb6e9cb),
	.w8(32'h3c54e78f),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5a4d1e),
	.w1(32'h3c9d6437),
	.w2(32'hbba99d83),
	.w3(32'h3bef0601),
	.w4(32'h3a8a9852),
	.w5(32'h3b22991c),
	.w6(32'h3b1eabd6),
	.w7(32'h3cca269c),
	.w8(32'hbb118989),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd6120f9),
	.w1(32'hba11c8fc),
	.w2(32'hbbb6a7a6),
	.w3(32'h3acc5b9d),
	.w4(32'h3914d0e6),
	.w5(32'h3bfb982b),
	.w6(32'hbc7b2496),
	.w7(32'hbab6c587),
	.w8(32'hbb5ad5cf),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf1f3f1),
	.w1(32'hbbb0467c),
	.w2(32'h3b79b422),
	.w3(32'h3b9bd0cc),
	.w4(32'h3c054a3d),
	.w5(32'hbd0d8946),
	.w6(32'hbd46b8a8),
	.w7(32'hbbb639ce),
	.w8(32'hbcaabf90),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b20da17),
	.w1(32'hbb23b995),
	.w2(32'hba2e5508),
	.w3(32'h3b2f3762),
	.w4(32'hbaf69122),
	.w5(32'h3b97ef08),
	.w6(32'h3b0faca6),
	.w7(32'h3ae58a87),
	.w8(32'hb94eedb1),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3c52c5),
	.w1(32'hbba34dab),
	.w2(32'hb94857fb),
	.w3(32'hbbafb342),
	.w4(32'h3cede9ed),
	.w5(32'hbb1cf3ee),
	.w6(32'h3cf8f47c),
	.w7(32'h3b93d151),
	.w8(32'h3c28274a),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbac40b8),
	.w1(32'hbbb7a1ab),
	.w2(32'h3b589450),
	.w3(32'hbc742d0d),
	.w4(32'hbb11dcb1),
	.w5(32'hbbad67c9),
	.w6(32'hba8c8481),
	.w7(32'hbbd04e17),
	.w8(32'hbaa51f3a),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7699af),
	.w1(32'hba7a70c6),
	.w2(32'hbb734b54),
	.w3(32'hbbe458b6),
	.w4(32'hbd2bb4ce),
	.w5(32'hbc139d97),
	.w6(32'hbaa50fe1),
	.w7(32'h3c0276e6),
	.w8(32'hba4819ea),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab77a3d),
	.w1(32'hbc57f831),
	.w2(32'hbb97aa9e),
	.w3(32'hbb1f1f6d),
	.w4(32'hbc14aa41),
	.w5(32'h3bc81b74),
	.w6(32'hbc9592db),
	.w7(32'hbbea5ddd),
	.w8(32'hbc6dbe87),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b37cf3a),
	.w1(32'h3b7c849d),
	.w2(32'hb9ba0778),
	.w3(32'h3a0966f1),
	.w4(32'h3b7ec224),
	.w5(32'h3a77299d),
	.w6(32'hb99eddb1),
	.w7(32'hba1108ff),
	.w8(32'h3c15770c),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0f5109),
	.w1(32'h3c524bfd),
	.w2(32'h3aeece7f),
	.w3(32'h3cabf8de),
	.w4(32'h3a2bd7e5),
	.w5(32'hbc0b9a1e),
	.w6(32'h3b814af9),
	.w7(32'h3c4fd429),
	.w8(32'h3bd2cb39),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule