module layer_10_featuremap_150(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb739a541),
	.w1(32'hb7b5dfd5),
	.w2(32'hb775e598),
	.w3(32'hb7cfccf3),
	.w4(32'hb7e3ca65),
	.w5(32'hb71f437f),
	.w6(32'hb846f88f),
	.w7(32'hb87697f8),
	.w8(32'hb7bcf46e),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb71d8d),
	.w1(32'hbba29d0b),
	.w2(32'hbaec78ac),
	.w3(32'hbb1b02dc),
	.w4(32'hbb0c3fd1),
	.w5(32'hb9bafd1d),
	.w6(32'h3a80016d),
	.w7(32'h3ac79891),
	.w8(32'h3b238ebd),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7202090),
	.w1(32'hb71606a4),
	.w2(32'hb7313dca),
	.w3(32'hb6fc20d7),
	.w4(32'hb6fda159),
	.w5(32'hb6a98dfb),
	.w6(32'hb781d37f),
	.w7(32'hb701e9d7),
	.w8(32'hb7887079),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ef536a),
	.w1(32'hba0bcff2),
	.w2(32'hb9831d7f),
	.w3(32'h392673cf),
	.w4(32'h396fd752),
	.w5(32'h39ad5779),
	.w6(32'hb9bf904d),
	.w7(32'hb82545d9),
	.w8(32'h39071a95),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb87a5561),
	.w1(32'hb817ada3),
	.w2(32'hb711303c),
	.w3(32'hb86c738f),
	.w4(32'hb82e03ed),
	.w5(32'hb438be3a),
	.w6(32'hb85d604c),
	.w7(32'hb8333673),
	.w8(32'hb72b28ff),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37d926b9),
	.w1(32'h36eca84a),
	.w2(32'h3697ba9f),
	.w3(32'hb645c51b),
	.w4(32'hb56962fa),
	.w5(32'hb69eab84),
	.w6(32'hb7b3074b),
	.w7(32'hb7a3db5d),
	.w8(32'hb7bed01e),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa05373),
	.w1(32'hbb20eeb1),
	.w2(32'hbb9f4340),
	.w3(32'hbb086b6c),
	.w4(32'hb81f8da2),
	.w5(32'h3adf8905),
	.w6(32'hbb078f77),
	.w7(32'h3a563b85),
	.w8(32'hb8dccfa3),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0d75a2),
	.w1(32'h3c776bfd),
	.w2(32'hbadaddb0),
	.w3(32'h3b84de56),
	.w4(32'h3b5a640f),
	.w5(32'h38ffecb9),
	.w6(32'h39e0e400),
	.w7(32'h3b6148a8),
	.w8(32'hbb0ca2a8),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad1ea72),
	.w1(32'h3a751a25),
	.w2(32'h39c10e2e),
	.w3(32'h3af25b0b),
	.w4(32'h3a0e23da),
	.w5(32'h390bdc47),
	.w6(32'h3b163b04),
	.w7(32'h39e82152),
	.w8(32'hba00ee61),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c14d5f7),
	.w1(32'h3b63de93),
	.w2(32'h3a3cd8a1),
	.w3(32'h3bde0ff0),
	.w4(32'h3aedf41c),
	.w5(32'h3b0d687f),
	.w6(32'h3b7f9f22),
	.w7(32'h3ac6db44),
	.w8(32'h3af0c3a2),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d14916),
	.w1(32'hb9e78dda),
	.w2(32'hb9806b89),
	.w3(32'hb981fd93),
	.w4(32'hba5e37aa),
	.w5(32'hba115c6b),
	.w6(32'h37f41d82),
	.w7(32'hba0f22b3),
	.w8(32'hb926ab09),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a90ede9),
	.w1(32'h3b24f15c),
	.w2(32'hbbd4967b),
	.w3(32'hbbd51947),
	.w4(32'hbb7c19a3),
	.w5(32'hbade8961),
	.w6(32'hbbbbefbd),
	.w7(32'hbb488b49),
	.w8(32'hbb878e32),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7bfe06),
	.w1(32'h3bcf5686),
	.w2(32'h3a436f23),
	.w3(32'h3c415266),
	.w4(32'h3bab644b),
	.w5(32'h39a02da6),
	.w6(32'h3aa40cd7),
	.w7(32'hbb1a8c15),
	.w8(32'hbbc551a3),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39aa2fbf),
	.w1(32'h3a43f53f),
	.w2(32'hba1295e8),
	.w3(32'h3a6bfd5b),
	.w4(32'h3aa0dbc5),
	.w5(32'h3af6a051),
	.w6(32'h3ae67369),
	.w7(32'h3a7301ad),
	.w8(32'h3b4d8d54),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb02c0c9),
	.w1(32'hba854ed2),
	.w2(32'h3a907259),
	.w3(32'h39d05f95),
	.w4(32'hba1158fc),
	.w5(32'h39ba9832),
	.w6(32'h3a94f555),
	.w7(32'h39dd941d),
	.w8(32'h3ab1804e),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba57448),
	.w1(32'hba8a3b6a),
	.w2(32'h3af4a219),
	.w3(32'h3b266715),
	.w4(32'h3b1284f4),
	.w5(32'h38310166),
	.w6(32'h3b77b4bf),
	.w7(32'h3a9c3ad7),
	.w8(32'h3accadca),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f95b7d),
	.w1(32'hb9caee13),
	.w2(32'hb9fb259c),
	.w3(32'h39aa7431),
	.w4(32'hba528c23),
	.w5(32'hba8647b9),
	.w6(32'h39dfe73d),
	.w7(32'hb99cc85d),
	.w8(32'hb9c92dbe),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c29a41e),
	.w1(32'h3bb93f6a),
	.w2(32'hbb35ecb4),
	.w3(32'h3b5cdef9),
	.w4(32'h3b286872),
	.w5(32'hb82c9c51),
	.w6(32'h3abd5966),
	.w7(32'hbb33daa7),
	.w8(32'hbbb3d7fa),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be42aaa),
	.w1(32'h3b6f8833),
	.w2(32'hbaaf0138),
	.w3(32'h3b973148),
	.w4(32'h3b323a62),
	.w5(32'hb9da1e52),
	.w6(32'h3a842004),
	.w7(32'hbaadd2d6),
	.w8(32'hbb77c490),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb854ac05),
	.w1(32'h389600fe),
	.w2(32'hb7afa4f6),
	.w3(32'h38add91e),
	.w4(32'hb8d1103a),
	.w5(32'hb81d574c),
	.w6(32'hb8c53752),
	.w7(32'hb919245f),
	.w8(32'hb805b0d4),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e377c0),
	.w1(32'h395deea5),
	.w2(32'h38c3af93),
	.w3(32'h37b2de1a),
	.w4(32'h390d9b99),
	.w5(32'h39013bd7),
	.w6(32'hb8a67eed),
	.w7(32'h3803b269),
	.w8(32'hb78f8a0b),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0368cc),
	.w1(32'hbacebdbe),
	.w2(32'h39553eee),
	.w3(32'hba5f8ff8),
	.w4(32'hba6bf66a),
	.w5(32'h38adfc52),
	.w6(32'hb99c496e),
	.w7(32'hb9d01c2e),
	.w8(32'h397a7474),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a88f635),
	.w1(32'h3bc08f17),
	.w2(32'h3c11e30b),
	.w3(32'hbb07d4f3),
	.w4(32'h3b35e271),
	.w5(32'hb9a9e132),
	.w6(32'hba4bd522),
	.w7(32'h3b700499),
	.w8(32'hba041e97),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af87d10),
	.w1(32'h390db695),
	.w2(32'h3ab9ef1d),
	.w3(32'h3b01d8e3),
	.w4(32'hb9efbf31),
	.w5(32'h3aeb4364),
	.w6(32'h3aa407be),
	.w7(32'hba45dea0),
	.w8(32'h3aaedba7),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc04b9fa),
	.w1(32'hbbeedf60),
	.w2(32'h3aea9cfb),
	.w3(32'hbadf3d03),
	.w4(32'hbba85941),
	.w5(32'h3ade1ec8),
	.w6(32'h3b96a0b6),
	.w7(32'h3abf4eda),
	.w8(32'h3b8e27af),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3949fc77),
	.w1(32'hb96d29f4),
	.w2(32'hb98dfd1e),
	.w3(32'h3a071700),
	.w4(32'hb91961bd),
	.w5(32'hb6a09f9b),
	.w6(32'h39258ccf),
	.w7(32'hb9c2b15f),
	.w8(32'h3912cbab),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ec0ca8),
	.w1(32'hb85d380d),
	.w2(32'hb899702f),
	.w3(32'hb8eae02c),
	.w4(32'hb86918ce),
	.w5(32'hb9194075),
	.w6(32'hb8fa60b2),
	.w7(32'hb8b8028c),
	.w8(32'hb91f4a7e),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aec2f1c),
	.w1(32'hbb74b218),
	.w2(32'hba2d8e12),
	.w3(32'h3b62fa40),
	.w4(32'h3b85e6a7),
	.w5(32'h3b4e036d),
	.w6(32'h3c149841),
	.w7(32'h3be9cca3),
	.w8(32'h3b25b711),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad0132f),
	.w1(32'hba82e5de),
	.w2(32'h3aa37b84),
	.w3(32'hbb45229d),
	.w4(32'hbb20ff98),
	.w5(32'hba6b8060),
	.w6(32'hbb35bb4b),
	.w7(32'hbb3329f0),
	.w8(32'hbaddf4b2),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb4597a),
	.w1(32'hbc1d0f4a),
	.w2(32'hbab47e87),
	.w3(32'h3b02cd41),
	.w4(32'hbacf17e6),
	.w5(32'h3bdaf011),
	.w6(32'h3bcaa833),
	.w7(32'h3b4eb626),
	.w8(32'h3bc84bb0),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6c42ef7),
	.w1(32'hb8ba3cc3),
	.w2(32'hb8a5588e),
	.w3(32'hb83ef6d6),
	.w4(32'hb908b8b6),
	.w5(32'hb8daafdb),
	.w6(32'hb7cd6dd8),
	.w7(32'hb8ab80bc),
	.w8(32'hb88a31fd),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h386b1842),
	.w1(32'hb746a9f9),
	.w2(32'hb85b4e9c),
	.w3(32'h36c68680),
	.w4(32'hb9220b21),
	.w5(32'hb9711a7a),
	.w6(32'h3931d536),
	.w7(32'hb8b23ed8),
	.w8(32'hb93a5c77),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab60aa1),
	.w1(32'h3a39cc98),
	.w2(32'hba558b4a),
	.w3(32'h3a2c30ef),
	.w4(32'hba30d81c),
	.w5(32'hba3f7874),
	.w6(32'hb91db0ff),
	.w7(32'hba97c1b2),
	.w8(32'hba6680cd),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4308b7),
	.w1(32'hbae77161),
	.w2(32'h395c12fd),
	.w3(32'hba045969),
	.w4(32'hba318b62),
	.w5(32'hb9326094),
	.w6(32'h39e312f1),
	.w7(32'h39bdb9e9),
	.w8(32'h3a8baadd),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39806162),
	.w1(32'hba07ad12),
	.w2(32'hba867b23),
	.w3(32'hb93e66e9),
	.w4(32'hb77d4611),
	.w5(32'hb98ef308),
	.w6(32'h3a38d567),
	.w7(32'h3a506bef),
	.w8(32'h37e6956e),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5fec94),
	.w1(32'h3b0e02fe),
	.w2(32'hb98ea185),
	.w3(32'h399f8453),
	.w4(32'h3a1f14de),
	.w5(32'h3a15632c),
	.w6(32'hba7e4cb1),
	.w7(32'hb8d6e2cc),
	.w8(32'hba91ff8d),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbabb08b),
	.w1(32'h3c7ec96f),
	.w2(32'hbbb6c364),
	.w3(32'hbc09c9bc),
	.w4(32'h3b1ee99e),
	.w5(32'hbba353d4),
	.w6(32'hbc0af48c),
	.w7(32'h3b7b38b1),
	.w8(32'hbb66683e),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe5c0cb),
	.w1(32'hbbedafcb),
	.w2(32'h3b1465a9),
	.w3(32'hbaedb2d3),
	.w4(32'hbbb3bc1b),
	.w5(32'hbaf88e9b),
	.w6(32'h3c018cfb),
	.w7(32'h3b0aba4b),
	.w8(32'h3b127edf),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc536d76),
	.w1(32'hbc47eb8d),
	.w2(32'h39b23a24),
	.w3(32'hbbd7b524),
	.w4(32'hbb9807be),
	.w5(32'h3ae07628),
	.w6(32'h3b4dce26),
	.w7(32'h3b584c8a),
	.w8(32'h3bc7465e),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bfe07c),
	.w1(32'h38f762d3),
	.w2(32'h3a9d625b),
	.w3(32'h3adfaadb),
	.w4(32'h3ad05178),
	.w5(32'h3abd8999),
	.w6(32'h3b1eaba5),
	.w7(32'h3b14225b),
	.w8(32'h3ad89571),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0d08fc),
	.w1(32'h39b50bde),
	.w2(32'h390443c6),
	.w3(32'h3a15f633),
	.w4(32'h398ba8aa),
	.w5(32'h391e749f),
	.w6(32'h39d06922),
	.w7(32'h39818316),
	.w8(32'h38913a84),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb86ba400),
	.w1(32'hb82b8596),
	.w2(32'hb83aebec),
	.w3(32'hb8a71bf0),
	.w4(32'hb829d86a),
	.w5(32'hb97ea873),
	.w6(32'hb8da7962),
	.w7(32'hb8d9fdc8),
	.w8(32'hb9b6463a),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba773be5),
	.w1(32'hbb21c850),
	.w2(32'hbb0d14ea),
	.w3(32'hbaa0ea4e),
	.w4(32'hbb36a014),
	.w5(32'hbb004578),
	.w6(32'hba86ae7f),
	.w7(32'hbb116511),
	.w8(32'hba657723),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3ee2a7),
	.w1(32'h3a326d85),
	.w2(32'h3ac0f6ea),
	.w3(32'h3bb98fab),
	.w4(32'h3ada1887),
	.w5(32'h390826d4),
	.w6(32'h3aeaefab),
	.w7(32'hbb615d8b),
	.w8(32'hbb18c822),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aae06ea),
	.w1(32'hba2ae587),
	.w2(32'h3b105d15),
	.w3(32'h3b438fb4),
	.w4(32'hba85a37a),
	.w5(32'h3a7a0e6a),
	.w6(32'h3b3838c0),
	.w7(32'hb9668189),
	.w8(32'h3a80e2b6),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad8fe08),
	.w1(32'h3b054508),
	.w2(32'h3adec19c),
	.w3(32'h3b3375a5),
	.w4(32'hba093996),
	.w5(32'h3a14ae9b),
	.w6(32'h3aaa2c46),
	.w7(32'hbaac2a46),
	.w8(32'hba06f342),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baf6a42),
	.w1(32'h3b23ba86),
	.w2(32'h3aff9fce),
	.w3(32'h3ba9359f),
	.w4(32'h3b05b3d6),
	.w5(32'h3a8fc407),
	.w6(32'h3bab69f0),
	.w7(32'h3b14316f),
	.w8(32'h3b117eca),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c819435),
	.w1(32'h3c159630),
	.w2(32'hba77b333),
	.w3(32'h3c2429d2),
	.w4(32'h3be62e97),
	.w5(32'h39e44213),
	.w6(32'h3984a757),
	.w7(32'h3aaa0cb0),
	.w8(32'hbbb46972),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94beaaf),
	.w1(32'hb9c8049a),
	.w2(32'h38909da8),
	.w3(32'hb9b08c7c),
	.w4(32'hba00c9c0),
	.w5(32'h39b471e9),
	.w6(32'hba1d4d9c),
	.w7(32'hb9a22fca),
	.w8(32'h3970efa1),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f39e24),
	.w1(32'hb903a0e7),
	.w2(32'h3a55d081),
	.w3(32'h38bd892c),
	.w4(32'h39ad9c96),
	.w5(32'h3aa7f71a),
	.w6(32'h39af5c1c),
	.w7(32'h39fb3b32),
	.w8(32'h3a83c98a),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa5f5d1),
	.w1(32'hba4d4a43),
	.w2(32'hb79bb0e7),
	.w3(32'hbae45592),
	.w4(32'hba9f19a2),
	.w5(32'h399371e1),
	.w6(32'hbaddb490),
	.w7(32'hba97ca99),
	.w8(32'hb91dfd3f),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6c1586),
	.w1(32'hbaded05f),
	.w2(32'h3aa207f0),
	.w3(32'h3ac45b48),
	.w4(32'h39ea9072),
	.w5(32'h39d95ba5),
	.w6(32'h3b07dd96),
	.w7(32'h39884a8b),
	.w8(32'hba2da19d),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92d9588),
	.w1(32'h3a50f8c5),
	.w2(32'h3a248b35),
	.w3(32'hbaac9a56),
	.w4(32'h395275ef),
	.w5(32'h3a25554a),
	.w6(32'hb9b243fb),
	.w7(32'h3a1aa97b),
	.w8(32'h3a12ac30),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c28133b),
	.w1(32'h3c042068),
	.w2(32'h3adaa5eb),
	.w3(32'h3bc3efe1),
	.w4(32'h3b7d9673),
	.w5(32'hb9ca9437),
	.w6(32'hbb224819),
	.w7(32'hbae797d6),
	.w8(32'hbb0afa35),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab34b1a),
	.w1(32'h3a15e2b8),
	.w2(32'h3a3a0684),
	.w3(32'hba287192),
	.w4(32'hbaa427e2),
	.w5(32'hba1dfc8a),
	.w6(32'hb8bf49d6),
	.w7(32'hbae74ce5),
	.w8(32'hbab73651),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0a10ea),
	.w1(32'hba203dd6),
	.w2(32'h3741ca78),
	.w3(32'hb8048224),
	.w4(32'hb9490e94),
	.w5(32'h399df14b),
	.w6(32'h385a44dd),
	.w7(32'h38bdb929),
	.w8(32'h3a1785ba),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7c0e6e5),
	.w1(32'h37cd3a77),
	.w2(32'h37bfcf53),
	.w3(32'hb7886754),
	.w4(32'hb65ac586),
	.w5(32'h37954486),
	.w6(32'hb7fb7b5c),
	.w7(32'hb50bca32),
	.w8(32'h3746f0cc),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e9197f),
	.w1(32'hb9a3c690),
	.w2(32'h386e3cf1),
	.w3(32'hb996cf0d),
	.w4(32'hb8ca3891),
	.w5(32'h380859c3),
	.w6(32'h39548a21),
	.w7(32'h395cacfd),
	.w8(32'h3991c358),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9da8b43),
	.w1(32'hba4efa0d),
	.w2(32'hba87a761),
	.w3(32'hba081fff),
	.w4(32'hba848108),
	.w5(32'hba9dd850),
	.w6(32'h3a022f12),
	.w7(32'hb9885f8d),
	.w8(32'hba0a5d7b),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5b0b6e),
	.w1(32'hba56accb),
	.w2(32'hba837713),
	.w3(32'h397ef6e5),
	.w4(32'hba2936db),
	.w5(32'hba4dec52),
	.w6(32'h3939f0fe),
	.w7(32'hb992cf7a),
	.w8(32'hba02c12d),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b557c0f),
	.w1(32'h39c7c14b),
	.w2(32'hbb0bb6ca),
	.w3(32'h3a856f3a),
	.w4(32'hba830e91),
	.w5(32'hbb1c434d),
	.w6(32'hbaa7bb0e),
	.w7(32'hbb15508f),
	.w8(32'hbb31b7f2),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b935202),
	.w1(32'hbb599146),
	.w2(32'h38ba519e),
	.w3(32'h3aef4b0c),
	.w4(32'h3a33631b),
	.w5(32'hbacf1748),
	.w6(32'h3bb32ba9),
	.w7(32'h39d88940),
	.w8(32'hbac8930d),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h382d2ecd),
	.w1(32'h3620aefa),
	.w2(32'h37416018),
	.w3(32'h380e2245),
	.w4(32'hb83a5cf3),
	.w5(32'hb848316b),
	.w6(32'hb81c3a11),
	.w7(32'hb874b66e),
	.w8(32'hb8cec2bb),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3791a3f5),
	.w1(32'h36da900e),
	.w2(32'hb715b8df),
	.w3(32'h38148058),
	.w4(32'h37a00653),
	.w5(32'hb69859d0),
	.w6(32'hb58e8139),
	.w7(32'hb6a32016),
	.w8(32'hb7eb59cf),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb954b914),
	.w1(32'hb930234e),
	.w2(32'hb7a87cfe),
	.w3(32'hb922f493),
	.w4(32'hb8a11696),
	.w5(32'h37e1fd1f),
	.w6(32'hb76fd5d1),
	.w7(32'hb8be2cee),
	.w8(32'h371ee54d),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6d8d8cc),
	.w1(32'h37c0aa54),
	.w2(32'hb88ef6cb),
	.w3(32'hb7ec1640),
	.w4(32'hb78c1fe7),
	.w5(32'hb8ce4307),
	.w6(32'hb8463171),
	.w7(32'hb88db353),
	.w8(32'hb9020443),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1cdd9e),
	.w1(32'h3ac7d60f),
	.w2(32'hbbcf2ea5),
	.w3(32'hbb1125ec),
	.w4(32'hba55a005),
	.w5(32'hbb728660),
	.w6(32'h3b621198),
	.w7(32'hba465869),
	.w8(32'hbaf164d6),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6bc546),
	.w1(32'h3ab8402f),
	.w2(32'h3b184270),
	.w3(32'hbba328a0),
	.w4(32'hba9d3aef),
	.w5(32'h3b01f48a),
	.w6(32'hba0c1c60),
	.w7(32'hbb456f7e),
	.w8(32'hbb00f9a2),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0cf120),
	.w1(32'hbafd3652),
	.w2(32'h398cf47c),
	.w3(32'hbb65afae),
	.w4(32'hbb702139),
	.w5(32'hbb202f77),
	.w6(32'h39a95830),
	.w7(32'hbb2bac13),
	.w8(32'hbb680eb9),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc14986c),
	.w1(32'hbc0c650e),
	.w2(32'h3b9c752f),
	.w3(32'hbb48789e),
	.w4(32'hbbc90566),
	.w5(32'h3b0c978e),
	.w6(32'h3bc33c49),
	.w7(32'h39df5983),
	.w8(32'h3ba3e30e),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36a3f8ff),
	.w1(32'h3810e368),
	.w2(32'hb85ffd07),
	.w3(32'hb75fb45f),
	.w4(32'hb5c4013f),
	.w5(32'hb887b08c),
	.w6(32'hb8842c46),
	.w7(32'hb8658d90),
	.w8(32'hb8c3ef75),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8814965),
	.w1(32'h36f86fb3),
	.w2(32'hb82fcfc2),
	.w3(32'hb7e8605a),
	.w4(32'h37ca06e8),
	.w5(32'hb87802dc),
	.w6(32'hb880c129),
	.w7(32'hb81946bd),
	.w8(32'hb8c74c65),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h387f2574),
	.w1(32'h38471694),
	.w2(32'hb886ec81),
	.w3(32'h385d4a80),
	.w4(32'h37f0f732),
	.w5(32'hb8c8cb59),
	.w6(32'hb804d1d7),
	.w7(32'hb85a1601),
	.w8(32'hb9070cf8),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1de811),
	.w1(32'h3ae6d0f2),
	.w2(32'hba8aae67),
	.w3(32'h3b3c402d),
	.w4(32'h3b0bba8c),
	.w5(32'hbabd8b4d),
	.w6(32'h3b0c8e79),
	.w7(32'h39a0451a),
	.w8(32'hbb45943d),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b41dd0),
	.w1(32'h3893d1ba),
	.w2(32'h3803a782),
	.w3(32'hb6b2447c),
	.w4(32'h3812a0d6),
	.w5(32'hb859ce11),
	.w6(32'hb8d5cc0c),
	.w7(32'hb72a4d58),
	.w8(32'hb8e5a929),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba40f6d),
	.w1(32'h3bceb632),
	.w2(32'hb9917096),
	.w3(32'h3b08b6ec),
	.w4(32'h3a07b93a),
	.w5(32'hba23cef6),
	.w6(32'hbafeb42e),
	.w7(32'hb9a05268),
	.w8(32'hbac61858),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3f15d5),
	.w1(32'h3c2ca3c6),
	.w2(32'h38f6af2e),
	.w3(32'h3a28787d),
	.w4(32'h3b719b5c),
	.w5(32'hbb127e95),
	.w6(32'h3997e280),
	.w7(32'hba327b3e),
	.w8(32'hbb914179),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd0486e),
	.w1(32'h3aaa3524),
	.w2(32'h3b21374c),
	.w3(32'h3bf866b8),
	.w4(32'h3b5bad6f),
	.w5(32'h3aa60b62),
	.w6(32'h3b48d629),
	.w7(32'h3a73f2b3),
	.w8(32'hbab2ed13),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae48b5e),
	.w1(32'h3a4a9a61),
	.w2(32'h3a5cc350),
	.w3(32'hb9250a00),
	.w4(32'hb8847a97),
	.w5(32'h3a9e5a29),
	.w6(32'hb9aa4040),
	.w7(32'hb95571d8),
	.w8(32'h3a9350b0),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbf29ee),
	.w1(32'h3b8e983e),
	.w2(32'hbb4fa892),
	.w3(32'hb9ec8c3b),
	.w4(32'hb99091be),
	.w5(32'hbaa9810d),
	.w6(32'h3b2a8197),
	.w7(32'h3b01dbcf),
	.w8(32'h3aef9a79),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b042d29),
	.w1(32'hbaa3da64),
	.w2(32'h3ab64c72),
	.w3(32'h3a6c0d1e),
	.w4(32'hba4ea3c9),
	.w5(32'hb9bd1407),
	.w6(32'h3b0979b7),
	.w7(32'hba08caa6),
	.w8(32'h39f10959),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b98f306),
	.w1(32'h3b165d85),
	.w2(32'hb961ae7f),
	.w3(32'h3b6ac2f3),
	.w4(32'h3afa93a1),
	.w5(32'h389903ed),
	.w6(32'h39b53ce2),
	.w7(32'hba105077),
	.w8(32'hbb0e6b5e),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb67b0aab),
	.w1(32'hb3f56592),
	.w2(32'h35f02cbb),
	.w3(32'h35402c68),
	.w4(32'hb525325e),
	.w5(32'h36efb410),
	.w6(32'hb63c623c),
	.w7(32'hb5ebf2dd),
	.w8(32'hb6a7d4c1),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb80abe91),
	.w1(32'hb7e5aa5f),
	.w2(32'h376a11eb),
	.w3(32'h37dce6fa),
	.w4(32'h3800c312),
	.w5(32'h379f6eca),
	.w6(32'h380e0dc3),
	.w7(32'h3851374a),
	.w8(32'h37cb1723),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37492863),
	.w1(32'hb79ee3ec),
	.w2(32'hb71d1306),
	.w3(32'h38000be2),
	.w4(32'h3488a560),
	.w5(32'hb58e5ed9),
	.w6(32'hb74360f4),
	.w7(32'hb72fe5f5),
	.w8(32'hb653a6fe),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4c306a),
	.w1(32'hb9a2fb07),
	.w2(32'h3928c26c),
	.w3(32'hb9738787),
	.w4(32'h399d7200),
	.w5(32'h39f64229),
	.w6(32'hb8fd6b78),
	.w7(32'h39ccbd35),
	.w8(32'h3a219ed8),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2b1f11),
	.w1(32'h39b79c8a),
	.w2(32'h3a4a50a0),
	.w3(32'hba77f6be),
	.w4(32'hbaa04d19),
	.w5(32'hbaebbd31),
	.w6(32'h3ac2a57f),
	.w7(32'h3a049094),
	.w8(32'h39cd17d9),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91aa18f),
	.w1(32'h399013bf),
	.w2(32'h37b0dd09),
	.w3(32'h389354ab),
	.w4(32'h3778b6d1),
	.w5(32'hb9b0281b),
	.w6(32'h3996881c),
	.w7(32'hb85c666d),
	.w8(32'hba06e834),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae57bec),
	.w1(32'hb9e80e32),
	.w2(32'h3aace008),
	.w3(32'hbad88026),
	.w4(32'hbae196e1),
	.w5(32'h394fc24d),
	.w6(32'hbac4134e),
	.w7(32'hbab9e7dd),
	.w8(32'h3a881239),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae1db43),
	.w1(32'h3b938c21),
	.w2(32'h3a82315b),
	.w3(32'hb8b6d3a0),
	.w4(32'h3a973f19),
	.w5(32'hbad5be1e),
	.w6(32'hbb8d693f),
	.w7(32'hbaaeccd4),
	.w8(32'hbb474cb9),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9cbf68),
	.w1(32'hbb598243),
	.w2(32'h3aecd9f0),
	.w3(32'hba6014bf),
	.w4(32'hba82dfb6),
	.w5(32'h3adf4760),
	.w6(32'h3aa4696f),
	.w7(32'h3a650e51),
	.w8(32'h3b037837),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c31c2d6),
	.w1(32'h3bb0e2a8),
	.w2(32'hbbd90111),
	.w3(32'hbb06144e),
	.w4(32'h39d3a6eb),
	.w5(32'hbbc8326f),
	.w6(32'hb9e73f4b),
	.w7(32'hba284666),
	.w8(32'hbb857a49),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaae97b5),
	.w1(32'h39511fbd),
	.w2(32'h3b0e9d09),
	.w3(32'hbaabd9e8),
	.w4(32'hba795838),
	.w5(32'h3a93741f),
	.w6(32'h3ae538cc),
	.w7(32'h3aac7a35),
	.w8(32'h3a4e3b89),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdbe2fe),
	.w1(32'h3b88332c),
	.w2(32'h3a7d5254),
	.w3(32'hbaeffc30),
	.w4(32'hba8d42a3),
	.w5(32'hba40aade),
	.w6(32'hbb153359),
	.w7(32'hbaee8107),
	.w8(32'h3a9416ab),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab0f862),
	.w1(32'hba9141ce),
	.w2(32'hba0da871),
	.w3(32'hbb068574),
	.w4(32'hb88cd230),
	.w5(32'h3918171f),
	.w6(32'h3ad38ffe),
	.w7(32'h3a3ee24b),
	.w8(32'h3b035246),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb35376f),
	.w1(32'hbb50bfe2),
	.w2(32'h3ab1228d),
	.w3(32'h3b849401),
	.w4(32'hb91b947f),
	.w5(32'h3b62803a),
	.w6(32'h3b89beae),
	.w7(32'h3b440ba4),
	.w8(32'h3b48a8d5),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5822b7),
	.w1(32'hba6fe5d0),
	.w2(32'hb7bc8701),
	.w3(32'hba483330),
	.w4(32'hba735f0c),
	.w5(32'h39eb5313),
	.w6(32'hba79b6b7),
	.w7(32'hba366865),
	.w8(32'hba2d0391),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b814b08),
	.w1(32'h3afde437),
	.w2(32'h3aaf5736),
	.w3(32'h3a7e305d),
	.w4(32'h3ad7b1fa),
	.w5(32'h3b351479),
	.w6(32'hba8ab1e8),
	.w7(32'hb90fba28),
	.w8(32'h38edf942),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1ec422),
	.w1(32'h3b83f6aa),
	.w2(32'hbba52331),
	.w3(32'hbb10f52b),
	.w4(32'hbb3cd147),
	.w5(32'hbbb4791c),
	.w6(32'h3a894add),
	.w7(32'hbaeb01d2),
	.w8(32'hbb9b0450),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc2afe9),
	.w1(32'h3c116776),
	.w2(32'h3c1dbe02),
	.w3(32'hbbb95aab),
	.w4(32'h3af5d79e),
	.w5(32'h3b0830c0),
	.w6(32'hb8e2be08),
	.w7(32'h3c1a73af),
	.w8(32'h3b2f73ab),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbfbf78),
	.w1(32'hbb83ae49),
	.w2(32'h3acb9a07),
	.w3(32'hbb1889af),
	.w4(32'hbb1cfbda),
	.w5(32'h3b4e7e36),
	.w6(32'h3c136cda),
	.w7(32'h3b8ae4fe),
	.w8(32'h3bf63e19),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7c93f9),
	.w1(32'hbb3578aa),
	.w2(32'h3b3d71e5),
	.w3(32'h3932d81c),
	.w4(32'hba91943c),
	.w5(32'h3b946c74),
	.w6(32'h3b02c4db),
	.w7(32'h3aedfe62),
	.w8(32'h3baa6f0c),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8f911f),
	.w1(32'h3bbe4bc0),
	.w2(32'hbc0548ca),
	.w3(32'hbc0fb5fc),
	.w4(32'hbbadb04b),
	.w5(32'hbb52ab33),
	.w6(32'hbbaaea8a),
	.w7(32'hbaf9c815),
	.w8(32'hbacc9b65),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3748dc6c),
	.w1(32'hba75f3c8),
	.w2(32'h39990aae),
	.w3(32'hb9b0bb25),
	.w4(32'hbb0e3184),
	.w5(32'hb8b44869),
	.w6(32'hba9dae11),
	.w7(32'hbb06a09d),
	.w8(32'hbab36ea0),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be85b33),
	.w1(32'h3c8b6ff2),
	.w2(32'h3b9063b4),
	.w3(32'h3b415c18),
	.w4(32'hbb529992),
	.w5(32'hba8c1da7),
	.w6(32'hbbf8ccf3),
	.w7(32'hbb0360a1),
	.w8(32'hbaf5260e),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4e7fb5),
	.w1(32'h3b8c4e32),
	.w2(32'hba5a7a65),
	.w3(32'hb8424e9d),
	.w4(32'hbac6e4c1),
	.w5(32'hb9d8a41f),
	.w6(32'h39b40c00),
	.w7(32'hbb267b64),
	.w8(32'hbadd731e),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb813dbc2),
	.w1(32'hb8374721),
	.w2(32'h38edfdf4),
	.w3(32'hb696c86a),
	.w4(32'hb88cb0e3),
	.w5(32'h38339573),
	.w6(32'h382232d8),
	.w7(32'hb8ca27e7),
	.w8(32'h38036d60),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6120da),
	.w1(32'hb9c00ded),
	.w2(32'h3a9c100f),
	.w3(32'hba22b7d3),
	.w4(32'hba0c60de),
	.w5(32'hb9f9a525),
	.w6(32'h3a9e57a4),
	.w7(32'h37cc1112),
	.w8(32'h3a1e9ecc),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baa5074),
	.w1(32'h3a7d742a),
	.w2(32'hba21c2f2),
	.w3(32'h3b750c9a),
	.w4(32'h3b108625),
	.w5(32'h3b01d16b),
	.w6(32'hba053abc),
	.w7(32'h39d41bb3),
	.w8(32'hba398899),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4f6de4),
	.w1(32'hbb66a189),
	.w2(32'h3b38b408),
	.w3(32'hba14b151),
	.w4(32'hbaa2d35f),
	.w5(32'h3b8396c4),
	.w6(32'h3a4bd679),
	.w7(32'h3ab4835e),
	.w8(32'h3b78ff99),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6af1f9),
	.w1(32'hba78b0ee),
	.w2(32'h3b1463f6),
	.w3(32'h3a6d011f),
	.w4(32'hb87e7c34),
	.w5(32'h3b0d6d1c),
	.w6(32'h3b206335),
	.w7(32'h3aaf0096),
	.w8(32'h3b20fbf4),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb77983d),
	.w1(32'hbb95b9e7),
	.w2(32'hbb226361),
	.w3(32'hbadab8ef),
	.w4(32'hbb244f17),
	.w5(32'hba88da8d),
	.w6(32'h3acd6e4f),
	.w7(32'h3ad0635d),
	.w8(32'h3b209e96),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c7bbde),
	.w1(32'h3b0ea2c9),
	.w2(32'hbb0929ff),
	.w3(32'h3b01be2f),
	.w4(32'hba7b0c64),
	.w5(32'hbb24ad71),
	.w6(32'hbaaea3b6),
	.w7(32'hbb290e2c),
	.w8(32'hbba6d865),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b98d7f1),
	.w1(32'h3aa5cd1b),
	.w2(32'h3a9448f7),
	.w3(32'h3b6761ce),
	.w4(32'h3b899fb0),
	.w5(32'h3ab17e35),
	.w6(32'h3b7b0775),
	.w7(32'h3b72f0f8),
	.w8(32'h3b8fe3f7),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3923990f),
	.w1(32'hba896c42),
	.w2(32'h39fabc7c),
	.w3(32'h39f6039b),
	.w4(32'hba4a448e),
	.w5(32'h3a6a7cea),
	.w6(32'hb8af8aac),
	.w7(32'hba15d1de),
	.w8(32'h3a8b4db5),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39837e01),
	.w1(32'h39326c82),
	.w2(32'h38bc4789),
	.w3(32'h39805103),
	.w4(32'h38d83728),
	.w5(32'hb7caa6dd),
	.w6(32'h393f4164),
	.w7(32'hb81008c1),
	.w8(32'h380901af),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9eab4f1),
	.w1(32'h389291fb),
	.w2(32'h37ac4841),
	.w3(32'h3870f58a),
	.w4(32'h39a507f4),
	.w5(32'hb9b1beff),
	.w6(32'h392e5369),
	.w7(32'h39859ce1),
	.w8(32'h3a157586),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb862a598),
	.w1(32'h38c3e1c1),
	.w2(32'h38ec0a2d),
	.w3(32'hb80e14a6),
	.w4(32'h37f5143a),
	.w5(32'h3832e5b0),
	.w6(32'hb67dc3a2),
	.w7(32'h369e9fdb),
	.w8(32'h38289e05),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38c8ce96),
	.w1(32'h389c0ed4),
	.w2(32'h382ea7fc),
	.w3(32'h385f6e24),
	.w4(32'h378c7152),
	.w5(32'h38a275d1),
	.w6(32'h3802934b),
	.w7(32'hb80c7ffe),
	.w8(32'hb8eabc16),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a91262a),
	.w1(32'hba9386e8),
	.w2(32'h399c7089),
	.w3(32'h3add35ba),
	.w4(32'hbadbcc5f),
	.w5(32'h38636e7b),
	.w6(32'h3a990d2d),
	.w7(32'hbaf5bcda),
	.w8(32'hb8794fdc),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395349ab),
	.w1(32'hb8848791),
	.w2(32'hb920327b),
	.w3(32'h39f7c38c),
	.w4(32'h3804e8fc),
	.w5(32'hb9334db6),
	.w6(32'h39a3dfb9),
	.w7(32'h3883c7c6),
	.w8(32'hb95c38a8),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc3775e),
	.w1(32'h3b8c4043),
	.w2(32'hba45f020),
	.w3(32'h3af961c3),
	.w4(32'h3ac85f08),
	.w5(32'h38586c2a),
	.w6(32'hba196023),
	.w7(32'hba228896),
	.w8(32'hbb009c2a),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba7c5a0),
	.w1(32'hbbd544ce),
	.w2(32'hbba1ca92),
	.w3(32'h3a914f2e),
	.w4(32'hbb16b7d6),
	.w5(32'hba502ecc),
	.w6(32'h3bd98866),
	.w7(32'h3b93acdd),
	.w8(32'h3b95f713),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91126e4),
	.w1(32'hb889f885),
	.w2(32'hb8a07dc0),
	.w3(32'hb827e8f2),
	.w4(32'hb734c888),
	.w5(32'hb81b76ee),
	.w6(32'hb7bf2e61),
	.w7(32'hb80c6974),
	.w8(32'hb867e741),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8edf69c),
	.w1(32'hb94f4b77),
	.w2(32'hb96d8f59),
	.w3(32'h38f318c6),
	.w4(32'hb80e00be),
	.w5(32'hb8939ad8),
	.w6(32'h38e2d3cb),
	.w7(32'h37abba88),
	.w8(32'hb8e1a978),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7bacbe3),
	.w1(32'hb8205949),
	.w2(32'hb7cb5b40),
	.w3(32'hb80023a9),
	.w4(32'hb87b0524),
	.w5(32'hb883e868),
	.w6(32'h363d9714),
	.w7(32'hb7f098bf),
	.w8(32'hb7a19c66),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4b6dd6),
	.w1(32'hbac1c8b3),
	.w2(32'h38dce883),
	.w3(32'h3a19242a),
	.w4(32'hb9050224),
	.w5(32'h3b004993),
	.w6(32'hba3c871a),
	.w7(32'h3a7e5b77),
	.w8(32'h3acba6e8),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb42c12d),
	.w1(32'h3a4543f8),
	.w2(32'hb9bb6036),
	.w3(32'h3aa9d6e3),
	.w4(32'h3b0185bc),
	.w5(32'h3be3a038),
	.w6(32'h3ab35d5c),
	.w7(32'hba92ddf4),
	.w8(32'hbb1e67dd),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1341a2),
	.w1(32'hba45f696),
	.w2(32'hba6aebd0),
	.w3(32'h3bedd88c),
	.w4(32'hbb3e7db5),
	.w5(32'hbab63ce9),
	.w6(32'hbbacdcf0),
	.w7(32'hbba2adc9),
	.w8(32'hbb49decd),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0f130b),
	.w1(32'hbb51949b),
	.w2(32'hbb7b5511),
	.w3(32'hba92f5dd),
	.w4(32'hbb30f522),
	.w5(32'hbb7030e5),
	.w6(32'hbb5a6c43),
	.w7(32'hbb7252b1),
	.w8(32'hbb53ac64),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb269ec1),
	.w1(32'h3a5b574e),
	.w2(32'hba7b05ad),
	.w3(32'hbb2f792a),
	.w4(32'hba4bcb07),
	.w5(32'hbaa0f20c),
	.w6(32'hb94c9870),
	.w7(32'hbac75fac),
	.w8(32'hbb208c81),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb10dedc),
	.w1(32'h39ca9b48),
	.w2(32'h3aac93c1),
	.w3(32'hbaa240c1),
	.w4(32'h3bb18cf0),
	.w5(32'h3bd6c14e),
	.w6(32'hbb50ec24),
	.w7(32'hbadca384),
	.w8(32'hba507cb2),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8d46a1),
	.w1(32'hbab946e6),
	.w2(32'h3b773ccd),
	.w3(32'h3c143c17),
	.w4(32'h399cd284),
	.w5(32'h3b3c14be),
	.w6(32'hbb38b890),
	.w7(32'hb9b4a6d8),
	.w8(32'hbad86607),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8fcf74),
	.w1(32'hbb977a18),
	.w2(32'h38f0bf5f),
	.w3(32'hbb81cc54),
	.w4(32'hbb80c012),
	.w5(32'h3a1e5e2e),
	.w6(32'hbb5ba6d6),
	.w7(32'h398855b6),
	.w8(32'h3a9b6e0c),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2b920e),
	.w1(32'h39986421),
	.w2(32'hbbd48a19),
	.w3(32'h3b91fb73),
	.w4(32'hbb31d751),
	.w5(32'hbbbe726a),
	.w6(32'hbb9544ab),
	.w7(32'hbbbc35cb),
	.w8(32'hbbda5b95),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc046b3b),
	.w1(32'hba85287b),
	.w2(32'h39f65b05),
	.w3(32'hbb98b194),
	.w4(32'h3a0a52b8),
	.w5(32'h3b9e87c5),
	.w6(32'h3b8f3a5b),
	.w7(32'h3b996fac),
	.w8(32'h3bf96f82),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c069b7c),
	.w1(32'h3b6179c9),
	.w2(32'h3ad2217f),
	.w3(32'h3bd17953),
	.w4(32'h3b739926),
	.w5(32'h3b0ef603),
	.w6(32'h3b1c60b5),
	.w7(32'h3b9d633b),
	.w8(32'h3afea9dc),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c37a358),
	.w1(32'hbb251c4d),
	.w2(32'hbbbe09c2),
	.w3(32'h3bbe4745),
	.w4(32'hbb931d6a),
	.w5(32'hbbe4e07a),
	.w6(32'hbbde97f4),
	.w7(32'hbc14adcb),
	.w8(32'hbc13c37b),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc38765b),
	.w1(32'hb9466b6f),
	.w2(32'h39281f19),
	.w3(32'hbc067d03),
	.w4(32'hbb7c2a92),
	.w5(32'hbb6293a4),
	.w6(32'hba8c5f46),
	.w7(32'hbb0dba8e),
	.w8(32'hbb69f39f),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9b4699),
	.w1(32'h3b97decc),
	.w2(32'h3b7280a3),
	.w3(32'hba6664e4),
	.w4(32'h3bb64937),
	.w5(32'h3c35daa8),
	.w6(32'hb96e8939),
	.w7(32'hba163724),
	.w8(32'h3b094445),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd77de2),
	.w1(32'hba95eb50),
	.w2(32'hb8d2bb32),
	.w3(32'h3c327d00),
	.w4(32'hbb0ee083),
	.w5(32'hbabd986c),
	.w6(32'hba9ab0e5),
	.w7(32'hba4e7841),
	.w8(32'hba1fda64),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb700df1),
	.w1(32'h3c07624e),
	.w2(32'h3c0ee30c),
	.w3(32'hb855da8a),
	.w4(32'h3c40cc37),
	.w5(32'h3c851bbb),
	.w6(32'h3c7bfd65),
	.w7(32'h3c88a57c),
	.w8(32'h3c880bde),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c65edf9),
	.w1(32'hbb3bfc00),
	.w2(32'hb9add73c),
	.w3(32'h3c60eb41),
	.w4(32'h363f6858),
	.w5(32'h3b760227),
	.w6(32'hbb493c6d),
	.w7(32'hbb665503),
	.w8(32'hbbd0f413),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae7decc),
	.w1(32'hb95c5408),
	.w2(32'h3a7e6b91),
	.w3(32'hb96dec6b),
	.w4(32'h3a5db15e),
	.w5(32'h3b60d220),
	.w6(32'hba0697c9),
	.w7(32'h3ab5a419),
	.w8(32'h3aaf26af),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5f4702),
	.w1(32'h3bc04a54),
	.w2(32'h3b40e3e3),
	.w3(32'h3b811b0a),
	.w4(32'h3b87da03),
	.w5(32'h3b397a5a),
	.w6(32'h3bb02e75),
	.w7(32'h3b75491a),
	.w8(32'h3b2d7016),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b85e7b4),
	.w1(32'h39f2d939),
	.w2(32'h39dee41d),
	.w3(32'h3aa934f5),
	.w4(32'h3a6a0b83),
	.w5(32'hba9d0d81),
	.w6(32'h38ada2a8),
	.w7(32'hbac79028),
	.w8(32'hbb06615f),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb779708),
	.w1(32'hba87fafe),
	.w2(32'hb984ee95),
	.w3(32'h39c145d8),
	.w4(32'hbaa7b310),
	.w5(32'hba52a646),
	.w6(32'h3ad43bc9),
	.w7(32'hba99b542),
	.w8(32'h393bb9ee),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be2d7da),
	.w1(32'h3bc4b0c9),
	.w2(32'h3ad9a243),
	.w3(32'h3be594be),
	.w4(32'h3be5b931),
	.w5(32'h3b93424b),
	.w6(32'h3b98d024),
	.w7(32'h3b42fa8d),
	.w8(32'hbb0af483),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6a9940),
	.w1(32'h3b532285),
	.w2(32'h3b33b42a),
	.w3(32'h3b8de4ff),
	.w4(32'h3b85a05a),
	.w5(32'h3bc9f09e),
	.w6(32'h3b4f6492),
	.w7(32'h3b6623a8),
	.w8(32'h3bcb8b9d),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c38aecd),
	.w1(32'h3b144dab),
	.w2(32'h3bb66062),
	.w3(32'h3c4f29db),
	.w4(32'h3b2ce01a),
	.w5(32'h3b8f734a),
	.w6(32'hbaeb4dcc),
	.w7(32'hbb68f047),
	.w8(32'hbb81b9ab),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b82bec7),
	.w1(32'hba96682f),
	.w2(32'hb99e5e43),
	.w3(32'h3aa90b6c),
	.w4(32'hb99d8d52),
	.w5(32'h3ad02b2f),
	.w6(32'hbad826c8),
	.w7(32'hba841a51),
	.w8(32'h3b1af731),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c370057),
	.w1(32'h3bec195f),
	.w2(32'hbb0815d9),
	.w3(32'h3b841815),
	.w4(32'h3b703aa0),
	.w5(32'h3a2fcb7e),
	.w6(32'h3a080467),
	.w7(32'h3a912daf),
	.w8(32'h3909e488),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbda707),
	.w1(32'hbc14264d),
	.w2(32'hbb0bf1db),
	.w3(32'h3be5a848),
	.w4(32'hbb2cea7a),
	.w5(32'hbba9f141),
	.w6(32'h3b41025a),
	.w7(32'hbb051f5c),
	.w8(32'hbba7ccc6),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc104df1),
	.w1(32'h3a068c90),
	.w2(32'hb9798ab4),
	.w3(32'hbbcde074),
	.w4(32'h3b16abee),
	.w5(32'h3b4a5da8),
	.w6(32'h3ae431ed),
	.w7(32'hbaf45abb),
	.w8(32'h3ab92a5b),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97f1742),
	.w1(32'hba80e26f),
	.w2(32'h37ba7bae),
	.w3(32'hbab58990),
	.w4(32'hbae54b3f),
	.w5(32'h3aebc288),
	.w6(32'hbac9403d),
	.w7(32'h372a86bf),
	.w8(32'h3b1dd600),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb9c8c0),
	.w1(32'hbb93cdd8),
	.w2(32'hbb7e6bcd),
	.w3(32'h3baed531),
	.w4(32'hbb946b9c),
	.w5(32'hbbae73db),
	.w6(32'hbb9bdfbc),
	.w7(32'hbbef0612),
	.w8(32'hbbe67fd3),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe7f67e),
	.w1(32'hbb97a124),
	.w2(32'hbb9ce2f4),
	.w3(32'hbba701a9),
	.w4(32'hbbbe3c99),
	.w5(32'hbbebafa2),
	.w6(32'hbba9eb61),
	.w7(32'hbbc76da1),
	.w8(32'hbb2bec12),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9f533b),
	.w1(32'hba4036d3),
	.w2(32'h39d5bb5d),
	.w3(32'hbb518503),
	.w4(32'h3abce0f3),
	.w5(32'h3a8eed04),
	.w6(32'h3b195255),
	.w7(32'h3ac87ffd),
	.w8(32'h3a8ab654),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae6e8c6),
	.w1(32'h3b6e3e2f),
	.w2(32'h3ace1d6b),
	.w3(32'h3a49d585),
	.w4(32'h3b22b9b8),
	.w5(32'h3b250c92),
	.w6(32'h3ac9b51b),
	.w7(32'h3aed70c4),
	.w8(32'h3b713403),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b574b48),
	.w1(32'hba241af3),
	.w2(32'hb8b9eea7),
	.w3(32'h3b6bb443),
	.w4(32'hba80b647),
	.w5(32'h3a0456e3),
	.w6(32'hba276e54),
	.w7(32'h39acd59f),
	.w8(32'h3b032ecb),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baff307),
	.w1(32'h3b9826bb),
	.w2(32'h3a763f4a),
	.w3(32'h3b315d46),
	.w4(32'h3b30795c),
	.w5(32'h3ab3efce),
	.w6(32'h3b505ddc),
	.w7(32'h3b8ba9cc),
	.w8(32'h3a1fd04b),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b08a858),
	.w1(32'hb9487e29),
	.w2(32'hbaaddb3f),
	.w3(32'h38a9b37b),
	.w4(32'hbb1c6b98),
	.w5(32'h39c93cb7),
	.w6(32'hba1302c5),
	.w7(32'hbb3b1377),
	.w8(32'hbbb83fc5),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b6a55),
	.w1(32'hbc20c14c),
	.w2(32'hbc146c2e),
	.w3(32'hb9881ed2),
	.w4(32'hbc100511),
	.w5(32'hbc13477b),
	.w6(32'hbb8b639d),
	.w7(32'hbc33499f),
	.w8(32'hbc37ede7),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc32a9d0),
	.w1(32'hbacbe280),
	.w2(32'hba2f918f),
	.w3(32'hbc078097),
	.w4(32'hbabaac53),
	.w5(32'hb928d0e3),
	.w6(32'hbb04927e),
	.w7(32'hbae5c079),
	.w8(32'hb8b461df),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6fd97f),
	.w1(32'hbc166933),
	.w2(32'hbb9ed6b8),
	.w3(32'hbb839c5b),
	.w4(32'hbbfc559e),
	.w5(32'hbbd32414),
	.w6(32'hbc1fc154),
	.w7(32'hbbb3b386),
	.w8(32'hbb901aed),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7a810a),
	.w1(32'hbb689401),
	.w2(32'hbb8054cb),
	.w3(32'hbb8c811c),
	.w4(32'hbb1d867f),
	.w5(32'hbb5f3f15),
	.w6(32'hbb01eee6),
	.w7(32'hbb83a36c),
	.w8(32'hbb5f31cb),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb917245),
	.w1(32'h3a3f1ec3),
	.w2(32'hba264f57),
	.w3(32'hbb5807f3),
	.w4(32'h3a492665),
	.w5(32'h3adc9b1e),
	.w6(32'h3a1a7d44),
	.w7(32'h3ace7c54),
	.w8(32'h3b2abdce),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b137bfe),
	.w1(32'hbba9b93e),
	.w2(32'hbb30a587),
	.w3(32'h3b44d7de),
	.w4(32'hbb9b79a8),
	.w5(32'hbb519b20),
	.w6(32'hbb2a2072),
	.w7(32'hbb758126),
	.w8(32'hbb250152),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb373598),
	.w1(32'h3b6b7cd2),
	.w2(32'hbb10e304),
	.w3(32'hbb641031),
	.w4(32'h3b1521a8),
	.w5(32'h39a1238f),
	.w6(32'h3a8947ec),
	.w7(32'h3a37f335),
	.w8(32'hb9032a11),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaec42de),
	.w1(32'hbb8da9f7),
	.w2(32'hbab8e80c),
	.w3(32'hbaec6e93),
	.w4(32'hbbe0e78f),
	.w5(32'hbbeeccf1),
	.w6(32'hbb935e87),
	.w7(32'hbb7a5d67),
	.w8(32'hbb8405f1),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbae9112),
	.w1(32'hbbeb5731),
	.w2(32'hbb391ad3),
	.w3(32'hbbbd47eb),
	.w4(32'hbb937084),
	.w5(32'h3a4ac38a),
	.w6(32'hb99c0dbf),
	.w7(32'hba68627e),
	.w8(32'h3b0f5a56),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a54d0fd),
	.w1(32'hbb8ed694),
	.w2(32'hbad1becf),
	.w3(32'hb89d5ea0),
	.w4(32'h3a935956),
	.w5(32'hbb3ed56f),
	.w6(32'h3a67b385),
	.w7(32'hbb38a2c4),
	.w8(32'hbb5f0a53),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd87861),
	.w1(32'h3b84e031),
	.w2(32'h3c11cf4f),
	.w3(32'h3ade83b3),
	.w4(32'h3b8ec59d),
	.w5(32'h3b3028f7),
	.w6(32'h3c0dacd6),
	.w7(32'h3b43661a),
	.w8(32'h39d34ff1),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c110ae0),
	.w1(32'h3957a55c),
	.w2(32'h3afb0187),
	.w3(32'h3b935ba6),
	.w4(32'hbb5d0128),
	.w5(32'hba63e087),
	.w6(32'hbb30c1a2),
	.w7(32'hbb65449c),
	.w8(32'hbb399659),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0524c9),
	.w1(32'hba64510a),
	.w2(32'h3aa813d2),
	.w3(32'hbb1a61f8),
	.w4(32'h3b35e5b2),
	.w5(32'h3bcd905e),
	.w6(32'hbb547421),
	.w7(32'hbb18ae45),
	.w8(32'hb9a24a60),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b211d2b),
	.w1(32'h3a3ff726),
	.w2(32'h39009456),
	.w3(32'h3b5d5d8c),
	.w4(32'hba63ba2e),
	.w5(32'hbaaffcea),
	.w6(32'h39a8dfa7),
	.w7(32'hba3da778),
	.w8(32'hbac364bd),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa523d0),
	.w1(32'h38e6b9b0),
	.w2(32'h3a1d522f),
	.w3(32'hba8e21fc),
	.w4(32'h3a76973d),
	.w5(32'h3b26a6cc),
	.w6(32'h3aecb961),
	.w7(32'h3b1bec25),
	.w8(32'h3b9736df),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3e71b6),
	.w1(32'h3b2c4392),
	.w2(32'h3a5adb20),
	.w3(32'h3b6bb0d5),
	.w4(32'h3b242e3a),
	.w5(32'h3b30aac4),
	.w6(32'h3b36476d),
	.w7(32'h3b542859),
	.w8(32'h3b81001a),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b524475),
	.w1(32'h3b362d50),
	.w2(32'h3b9e8b5b),
	.w3(32'h3b517c44),
	.w4(32'h3b90afb7),
	.w5(32'h3bb5519e),
	.w6(32'hb9458f96),
	.w7(32'hb9fcda14),
	.w8(32'hbb2adf16),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91ee8fa),
	.w1(32'hbb605672),
	.w2(32'hbaf05480),
	.w3(32'h3a3bddfc),
	.w4(32'hba81765a),
	.w5(32'h3b5989ea),
	.w6(32'hbb94f13b),
	.w7(32'hbb241c50),
	.w8(32'hba758e54),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5270e0),
	.w1(32'hbb57bd19),
	.w2(32'hbafc5c1d),
	.w3(32'h3c55acb2),
	.w4(32'h39302380),
	.w5(32'h39d550e5),
	.w6(32'hbb67e635),
	.w7(32'hbad3096f),
	.w8(32'hba88dfc8),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba92f28b),
	.w1(32'hbc2788b4),
	.w2(32'hbb965645),
	.w3(32'h3a764299),
	.w4(32'hbc2456ee),
	.w5(32'hbbb5035e),
	.w6(32'hbc17b4ed),
	.w7(32'hbbd49994),
	.w8(32'hbbd0af8f),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f4c9d),
	.w1(32'hba98e0a1),
	.w2(32'hbb143127),
	.w3(32'hbbb2c50d),
	.w4(32'hba928957),
	.w5(32'hbb04f5de),
	.w6(32'hba938e99),
	.w7(32'hbb34f1ef),
	.w8(32'hbb22a87d),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6bd6b0),
	.w1(32'hbb3f485a),
	.w2(32'hbad04f1c),
	.w3(32'hbb0a1cc2),
	.w4(32'hbb0c9de4),
	.w5(32'hbb3a59ff),
	.w6(32'h3a095a4d),
	.w7(32'hbb505ffb),
	.w8(32'hba47237e),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8597c5),
	.w1(32'hb9fc77fc),
	.w2(32'hbb5701f0),
	.w3(32'hbb7dbf7d),
	.w4(32'hbba3a03a),
	.w5(32'hbb896379),
	.w6(32'hbbf60047),
	.w7(32'hbbbb2bf0),
	.w8(32'hbbdb48bc),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a1a0a),
	.w1(32'h3c39898f),
	.w2(32'h3c01fa6a),
	.w3(32'hbaec302d),
	.w4(32'h3be32575),
	.w5(32'h3c1b5956),
	.w6(32'h38525b91),
	.w7(32'h3b44ef3f),
	.w8(32'hbb116e03),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3a6d7f),
	.w1(32'hbbaaced9),
	.w2(32'hbba93c86),
	.w3(32'hbb02ca4d),
	.w4(32'hbb8a2875),
	.w5(32'hbb96ee55),
	.w6(32'hbb9fb67c),
	.w7(32'hbbc75bcb),
	.w8(32'hbbb6a35c),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c654e20),
	.w1(32'h3c1295ee),
	.w2(32'hbb04aae0),
	.w3(32'h3c00ea94),
	.w4(32'h3a5926a4),
	.w5(32'hbbb28d71),
	.w6(32'hbb0934c9),
	.w7(32'hbc63966c),
	.w8(32'hbc8f7996),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf3a67f),
	.w1(32'hbc10a070),
	.w2(32'hbbb324a3),
	.w3(32'h3b8eb0f7),
	.w4(32'hbba62252),
	.w5(32'hbc233f81),
	.w6(32'h3ba72f3b),
	.w7(32'hbaf0c805),
	.w8(32'hbbb42ec6),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8cb42b),
	.w1(32'h3b5e67df),
	.w2(32'h391a688a),
	.w3(32'hbb9e5348),
	.w4(32'hbab235c4),
	.w5(32'hbb0f1caf),
	.w6(32'h3ab2b440),
	.w7(32'h3b7dc2e8),
	.w8(32'h3bada0c5),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb9556b),
	.w1(32'h3b127615),
	.w2(32'h3bdc708a),
	.w3(32'h3b057ab2),
	.w4(32'h3b35e9fa),
	.w5(32'h3bb9f78d),
	.w6(32'h3b0719bb),
	.w7(32'h3bc04a53),
	.w8(32'h3a1c017f),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2d21de),
	.w1(32'hbb6f2830),
	.w2(32'hbb1fc130),
	.w3(32'h3b117cef),
	.w4(32'hbaba744e),
	.w5(32'hbb39e071),
	.w6(32'hbac2b3bc),
	.w7(32'hbb735173),
	.w8(32'hbb73ba53),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbeefc0),
	.w1(32'hbade185c),
	.w2(32'hba976787),
	.w3(32'hbb889c30),
	.w4(32'hba50ebea),
	.w5(32'hba64b479),
	.w6(32'hba8863c7),
	.w7(32'hba7bd050),
	.w8(32'hba35c151),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb015475),
	.w1(32'h3b822def),
	.w2(32'h3b1ffc97),
	.w3(32'hbb3acf98),
	.w4(32'h3b32a6ea),
	.w5(32'h3ba18a40),
	.w6(32'hba5b50d5),
	.w7(32'h3b46721b),
	.w8(32'hba4a486c),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb797296),
	.w1(32'h3b86063c),
	.w2(32'h3b184d91),
	.w3(32'hbbd17d07),
	.w4(32'h3b13de10),
	.w5(32'h39b41463),
	.w6(32'h3b431dc1),
	.w7(32'h3b4ae5e2),
	.w8(32'h3ae98140),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7f881a),
	.w1(32'hba03ddf4),
	.w2(32'hb9a9f490),
	.w3(32'h3ba524f5),
	.w4(32'h3a7fa920),
	.w5(32'hb9ea25ae),
	.w6(32'h3b7ae4ef),
	.w7(32'h398d342c),
	.w8(32'hb7ca21aa),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad52d3d),
	.w1(32'h3a9cf626),
	.w2(32'h3a689091),
	.w3(32'hbaf6a6f0),
	.w4(32'h39fde3f9),
	.w5(32'h3b5b7515),
	.w6(32'h3985cdf7),
	.w7(32'h3a8194b0),
	.w8(32'h3b3bdb5f),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c43b450),
	.w1(32'h3bf56460),
	.w2(32'h3bca0509),
	.w3(32'h3c1cfe6c),
	.w4(32'h3c054d40),
	.w5(32'h3bd310cb),
	.w6(32'hba315c0b),
	.w7(32'hbabcc9e4),
	.w8(32'hbbc65aac),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3d916d),
	.w1(32'h3abdc5c1),
	.w2(32'hb9a2ecec),
	.w3(32'hbb866dfa),
	.w4(32'hbad8fe4f),
	.w5(32'hbb1aba62),
	.w6(32'hb9b44928),
	.w7(32'hbb313f00),
	.w8(32'hbb60d8a8),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9dc85b),
	.w1(32'hb90c05a2),
	.w2(32'hba2f25f5),
	.w3(32'hbb2eb69b),
	.w4(32'hb928cc59),
	.w5(32'h3a9a3b5d),
	.w6(32'hb914e070),
	.w7(32'h3a560f0b),
	.w8(32'h3b1436a8),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b849e31),
	.w1(32'h3b27b2c6),
	.w2(32'hbaabe3ee),
	.w3(32'h3b7cf19d),
	.w4(32'h37f109ba),
	.w5(32'h3ad34dca),
	.w6(32'h384ba13c),
	.w7(32'h38b867e6),
	.w8(32'h3b37b919),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b093519),
	.w1(32'h3a62fc4a),
	.w2(32'h398bba55),
	.w3(32'h3b1edde6),
	.w4(32'h3a2852a6),
	.w5(32'h3b0f7405),
	.w6(32'h39abe617),
	.w7(32'h3a306bc5),
	.w8(32'h3b2d876f),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bca02e7),
	.w1(32'hbb94fcbe),
	.w2(32'hbbf27ee4),
	.w3(32'h3bdd8ec9),
	.w4(32'hbbce7c5a),
	.w5(32'hbc15ae84),
	.w6(32'hbbb7c280),
	.w7(32'hbbee6459),
	.w8(32'hbc0eb187),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc32de27),
	.w1(32'hbbd89780),
	.w2(32'hba9d1f68),
	.w3(32'hbc0197d8),
	.w4(32'hbb8289c7),
	.w5(32'hbadd8cce),
	.w6(32'hbb5a1aa3),
	.w7(32'hbbef0b61),
	.w8(32'hbbaa8319),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a54b627),
	.w1(32'h3b6698c6),
	.w2(32'h3b4b77f5),
	.w3(32'h3ad5f4aa),
	.w4(32'h3b81b5af),
	.w5(32'h3bae0940),
	.w6(32'h3ba19ac6),
	.w7(32'h3ba0b900),
	.w8(32'h3bdff96c),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb2160b),
	.w1(32'hbb3a2e13),
	.w2(32'hbb5f3c6c),
	.w3(32'h3ba12ed6),
	.w4(32'hbb309329),
	.w5(32'hbb7c4d08),
	.w6(32'hbb2c6db6),
	.w7(32'hbb91f625),
	.w8(32'hbbc05b84),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc15e36b),
	.w1(32'hbaaf2227),
	.w2(32'hbacb5c26),
	.w3(32'hbbb6b93a),
	.w4(32'h3a6f30b2),
	.w5(32'h3ae77f3c),
	.w6(32'h3b997aca),
	.w7(32'hb88c3244),
	.w8(32'h3b1a1210),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba39b6f),
	.w1(32'h3b8c235c),
	.w2(32'h3b367921),
	.w3(32'h3b9428c3),
	.w4(32'h3b9fb929),
	.w5(32'h3bce998b),
	.w6(32'h3b5073b2),
	.w7(32'h3b9026a9),
	.w8(32'h3bbb74a6),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c901d17),
	.w1(32'h3b8cf480),
	.w2(32'hbae1b9ef),
	.w3(32'h3c93dba1),
	.w4(32'h3b82610b),
	.w5(32'hbb7eaaf1),
	.w6(32'h3b83aac7),
	.w7(32'hbb5fbd56),
	.w8(32'hbb8275c9),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad77906),
	.w1(32'hbb89ae09),
	.w2(32'hbb2a39ad),
	.w3(32'hbab27985),
	.w4(32'hbb9757dd),
	.w5(32'hbb5dfd98),
	.w6(32'hbb9edc74),
	.w7(32'hbb858ad6),
	.w8(32'hbb8b4a2a),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb725ccd),
	.w1(32'hbae0eaa0),
	.w2(32'hbaca42f7),
	.w3(32'hbb760254),
	.w4(32'hbb265ec6),
	.w5(32'hbb32b1a0),
	.w6(32'hbb56e72f),
	.w7(32'hbb4b6229),
	.w8(32'hbb7e0cc5),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb65ed15),
	.w1(32'hba54c380),
	.w2(32'hbbc45a05),
	.w3(32'hbbb00a23),
	.w4(32'hbbc0a340),
	.w5(32'hbc066c34),
	.w6(32'hbba6ce95),
	.w7(32'hbc07ece9),
	.w8(32'hbc2c965a),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcffef3),
	.w1(32'h3b82d663),
	.w2(32'h3b5cfc81),
	.w3(32'hbbff6fcb),
	.w4(32'hbaaaea14),
	.w5(32'hb9bd2180),
	.w6(32'h3b0273f3),
	.w7(32'h3a9c34e4),
	.w8(32'h3a866804),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a86e15c),
	.w1(32'h3b622015),
	.w2(32'h3b92846c),
	.w3(32'hb915708c),
	.w4(32'h3b60cb50),
	.w5(32'h3b6afe3b),
	.w6(32'h3b9959f8),
	.w7(32'h3b428938),
	.w8(32'h3b34a52c),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1a8c98),
	.w1(32'hba3dd42f),
	.w2(32'hbc0b0718),
	.w3(32'hbbad6e0d),
	.w4(32'hbc07133c),
	.w5(32'hbb94ae8c),
	.w6(32'hbc085628),
	.w7(32'hbc015832),
	.w8(32'hbc0093ed),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb642685),
	.w1(32'h3ab1a1c5),
	.w2(32'h3aeaa822),
	.w3(32'hba30cd0b),
	.w4(32'h3b2152a5),
	.w5(32'h3b74bfc4),
	.w6(32'h3b2e9fe3),
	.w7(32'h3b27f068),
	.w8(32'h3b83d3ef),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8eb9f6),
	.w1(32'hbaf97531),
	.w2(32'hbb871709),
	.w3(32'h3bb5012a),
	.w4(32'hbb2bd769),
	.w5(32'hbb58be3e),
	.w6(32'hbb27e9ba),
	.w7(32'hbb5dcabc),
	.w8(32'hbb774a0f),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0fa1f5),
	.w1(32'h3bc0ba46),
	.w2(32'h389dacd5),
	.w3(32'hbc1a49b8),
	.w4(32'h3b446d55),
	.w5(32'h3b51c01c),
	.w6(32'hbb86b69d),
	.w7(32'h3b27ddf8),
	.w8(32'h3b8c1b6c),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca598e5),
	.w1(32'h3c102355),
	.w2(32'h399450b7),
	.w3(32'h3c87f192),
	.w4(32'h3b195bcb),
	.w5(32'hbb9c295c),
	.w6(32'h38d8ee1c),
	.w7(32'hbb9289f4),
	.w8(32'hbc0b6fc1),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be5fe05),
	.w1(32'h3bd09bf8),
	.w2(32'h39aeb23b),
	.w3(32'h3a302ef1),
	.w4(32'h3b5f3d89),
	.w5(32'h3b1177db),
	.w6(32'h3a3b6eb0),
	.w7(32'h3b178a13),
	.w8(32'h3b051fdd),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba564e1b),
	.w1(32'hbbed3fd7),
	.w2(32'hbb8fbad5),
	.w3(32'h3a947378),
	.w4(32'hbb9ef3e9),
	.w5(32'hbb54c2fc),
	.w6(32'hbab4be8b),
	.w7(32'hbb7a8900),
	.w8(32'hbb9887de),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0be5cf),
	.w1(32'hbbf54553),
	.w2(32'hbb582f0f),
	.w3(32'hbb9b91ed),
	.w4(32'hbbca5ebc),
	.w5(32'hbba31a4b),
	.w6(32'hba902ef7),
	.w7(32'hbb8ae35f),
	.w8(32'hba3e1085),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb17d32e),
	.w1(32'hbb297bbc),
	.w2(32'hbb033fe1),
	.w3(32'hbade0678),
	.w4(32'hbac1a58e),
	.w5(32'hbaa98b93),
	.w6(32'hbad75b8e),
	.w7(32'hbb083784),
	.w8(32'hbb0be1d4),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb113b87),
	.w1(32'hbba3cbf1),
	.w2(32'h3a3d5624),
	.w3(32'hba682c80),
	.w4(32'hbc030f5c),
	.w5(32'hbb3347c6),
	.w6(32'hbbeba9de),
	.w7(32'hbb3b6056),
	.w8(32'hbb6d11f4),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb991f16a),
	.w1(32'h387e87bf),
	.w2(32'hbaa1dd8c),
	.w3(32'hbb5d0fdd),
	.w4(32'h3b2638de),
	.w5(32'h3a943e2b),
	.w6(32'h3ad0e097),
	.w7(32'h3a266930),
	.w8(32'hba54acd9),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a576d05),
	.w1(32'h3aa07f64),
	.w2(32'h3a2f767f),
	.w3(32'h3ad1ee67),
	.w4(32'h3b1b8042),
	.w5(32'h3afa85d5),
	.w6(32'h3a065841),
	.w7(32'h3a061dad),
	.w8(32'hbb00892f),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4f6f0d),
	.w1(32'hbbac96ab),
	.w2(32'hbbad1038),
	.w3(32'h3a16a22e),
	.w4(32'hbb9d41ac),
	.w5(32'hbb955f06),
	.w6(32'hbbabc507),
	.w7(32'hbb846636),
	.w8(32'hbb8fc553),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaec7ff),
	.w1(32'hbbdf0467),
	.w2(32'hbb8fb91c),
	.w3(32'hbbd4ed90),
	.w4(32'hbbe4cd56),
	.w5(32'hbb94264c),
	.w6(32'hbc04a1ed),
	.w7(32'hbbd218fd),
	.w8(32'hbc185d04),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc012ec8),
	.w1(32'hbafbf0d6),
	.w2(32'h3bbc9010),
	.w3(32'hbbca1604),
	.w4(32'hba86428c),
	.w5(32'h3b9f3c1b),
	.w6(32'hba8dee0c),
	.w7(32'h3a97a492),
	.w8(32'hbb0d1cd3),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3710feb0),
	.w1(32'hbb2345e4),
	.w2(32'h3ba11def),
	.w3(32'hba63e59d),
	.w4(32'hbb8d3280),
	.w5(32'h3aa8ed70),
	.w6(32'hba81a671),
	.w7(32'h3afffce5),
	.w8(32'hb9cce492),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c403057),
	.w1(32'h3c6ca51e),
	.w2(32'h39d3fa0d),
	.w3(32'hbaee00fb),
	.w4(32'h3c2343a6),
	.w5(32'h3c01a183),
	.w6(32'h3bed4050),
	.w7(32'h3c167091),
	.w8(32'h3baf7639),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c335326),
	.w1(32'h3b23c004),
	.w2(32'h3986378f),
	.w3(32'h3c119c83),
	.w4(32'h3abf34ba),
	.w5(32'h3b1e76a3),
	.w6(32'h3a923ba1),
	.w7(32'h3b36d54a),
	.w8(32'h3b4a4dbd),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2ac6c5),
	.w1(32'h3b434215),
	.w2(32'h3ab5f21d),
	.w3(32'h3b605110),
	.w4(32'h3b4a87f1),
	.w5(32'h3b525241),
	.w6(32'h3b40c690),
	.w7(32'h3b5c5fa2),
	.w8(32'h3b808d44),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3912e4),
	.w1(32'h3b86a40c),
	.w2(32'hba75781b),
	.w3(32'h3bdba4f7),
	.w4(32'h3b07bca3),
	.w5(32'h3b074477),
	.w6(32'h3ac84494),
	.w7(32'h3aeafec1),
	.w8(32'h3a8d0cac),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b14b3c9),
	.w1(32'hbb6b7073),
	.w2(32'hbb41a173),
	.w3(32'h3b44e6d5),
	.w4(32'hbb2aefea),
	.w5(32'hbb1bef0e),
	.w6(32'hbb312ba2),
	.w7(32'hbb22d6dc),
	.w8(32'hbb07d0f6),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5c039a),
	.w1(32'h3b93e436),
	.w2(32'h3b62d5ab),
	.w3(32'hbb3ba071),
	.w4(32'h3b80e7bc),
	.w5(32'h3b92cceb),
	.w6(32'h3b57ea8d),
	.w7(32'h3b3bc7b7),
	.w8(32'h3ba6b384),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be91419),
	.w1(32'h3b785528),
	.w2(32'h3b0eafb0),
	.w3(32'h3bfbafb2),
	.w4(32'h3b74dd00),
	.w5(32'h3b77d746),
	.w6(32'h3b6c019f),
	.w7(32'h3b88d147),
	.w8(32'h3b9a30d1),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b93805f),
	.w1(32'hbbc5ff96),
	.w2(32'h37c5cd5b),
	.w3(32'h3b83246e),
	.w4(32'hbba6c77d),
	.w5(32'hbae53ff0),
	.w6(32'hbbc6b91b),
	.w7(32'hbb6ef301),
	.w8(32'hbb443c49),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9061ef),
	.w1(32'hbab26fdd),
	.w2(32'hb98aa355),
	.w3(32'hb97d9faf),
	.w4(32'h39e27682),
	.w5(32'h3b31fbb4),
	.w6(32'h3a4f6277),
	.w7(32'h3aa19e4a),
	.w8(32'h3afe7b71),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4cda5d),
	.w1(32'hbb2451f6),
	.w2(32'h3ba3bc8b),
	.w3(32'h3bf608fc),
	.w4(32'hb8c810c5),
	.w5(32'h3b303885),
	.w6(32'hb978f4b6),
	.w7(32'h394c91c3),
	.w8(32'h3b212c59),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c791ad8),
	.w1(32'h3ace2eb4),
	.w2(32'hb94b0dc6),
	.w3(32'h3bfddbb1),
	.w4(32'hba9fef03),
	.w5(32'h3b18cccc),
	.w6(32'hbb7e2dee),
	.w7(32'hbb06abaa),
	.w8(32'h3764856f),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5047a0),
	.w1(32'hbabd33e0),
	.w2(32'hbbc2a24b),
	.w3(32'h3bff954c),
	.w4(32'hbaf76588),
	.w5(32'hbc03d56d),
	.w6(32'hbbb6b0d6),
	.w7(32'hbbde5cb4),
	.w8(32'hbc16dd34),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd71437),
	.w1(32'hbb86bbb3),
	.w2(32'hbac8e032),
	.w3(32'hbbb3e93a),
	.w4(32'hbb67da4c),
	.w5(32'hba41d91e),
	.w6(32'hbb585053),
	.w7(32'hbaffe5c5),
	.w8(32'hba08887c),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b38f4f5),
	.w1(32'h3b9e4306),
	.w2(32'h3b1e159f),
	.w3(32'h3acaa833),
	.w4(32'h3bb51984),
	.w5(32'h3bb18fd7),
	.w6(32'h3ba0e654),
	.w7(32'h3bc3fc56),
	.w8(32'h3bdc0b4a),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcdb47c),
	.w1(32'h3aaf497e),
	.w2(32'hb9b084a1),
	.w3(32'h3bbdf774),
	.w4(32'h3a600d8c),
	.w5(32'h3a8e469b),
	.w6(32'h3adbc4cf),
	.w7(32'h3b1110be),
	.w8(32'h3b32402a),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b04f6fb),
	.w1(32'h3ae203da),
	.w2(32'h39ecf416),
	.w3(32'h3b027cb8),
	.w4(32'h3aafa265),
	.w5(32'h3b00cbb2),
	.w6(32'h3b03d2a6),
	.w7(32'h3b35e477),
	.w8(32'h3b4a3c6b),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba62a36),
	.w1(32'h3b845500),
	.w2(32'h3c24fb7d),
	.w3(32'h3b7137f7),
	.w4(32'h391fabb3),
	.w5(32'h3a900680),
	.w6(32'h3b628889),
	.w7(32'h3bd28b75),
	.w8(32'h3bb76b67),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1c45b0),
	.w1(32'hba04e10c),
	.w2(32'h3973e717),
	.w3(32'h3901de03),
	.w4(32'h3a8554cd),
	.w5(32'h3a460c23),
	.w6(32'h3aebf055),
	.w7(32'hba3b8eec),
	.w8(32'h38c553fe),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a5bd9c),
	.w1(32'hbc2106b7),
	.w2(32'hbc002144),
	.w3(32'hb95fb0db),
	.w4(32'hbc1f1f9c),
	.w5(32'hbbd99168),
	.w6(32'hbc2d79b9),
	.w7(32'hbc11d8b3),
	.w8(32'hbbef9c65),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc69e0f),
	.w1(32'hbb94978d),
	.w2(32'hbb5564e0),
	.w3(32'hbb958a0d),
	.w4(32'hbb9d1252),
	.w5(32'hbb4684f4),
	.w6(32'hbbb13ad4),
	.w7(32'hbb89f4a2),
	.w8(32'hbb9309b5),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6e920b),
	.w1(32'h3ae70148),
	.w2(32'hb93bc968),
	.w3(32'hbad25754),
	.w4(32'h3b009928),
	.w5(32'h3b129a73),
	.w6(32'h3b04013d),
	.w7(32'h3b276f22),
	.w8(32'h3b539129),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbb866b),
	.w1(32'hb781be88),
	.w2(32'h3bcd6267),
	.w3(32'h3bb5e1e4),
	.w4(32'hbb0dcf82),
	.w5(32'h3a9de47c),
	.w6(32'hb9dfaba1),
	.w7(32'h3b2c4f3f),
	.w8(32'hb983201f),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b341901),
	.w1(32'hbc18d4a5),
	.w2(32'hbbb35965),
	.w3(32'hbb0d371e),
	.w4(32'hbc172422),
	.w5(32'hbb8fe70e),
	.w6(32'hbc42bfe1),
	.w7(32'hbbedb86f),
	.w8(32'hbbf767d9),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b61f43a),
	.w1(32'hba9b6be2),
	.w2(32'hb98cf66f),
	.w3(32'hbb17d9bb),
	.w4(32'h3b22d2b4),
	.w5(32'hbb18ac48),
	.w6(32'h3b3775e7),
	.w7(32'hb9f62d2a),
	.w8(32'hba531391),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a83a581),
	.w1(32'h3949b55c),
	.w2(32'h370e80ec),
	.w3(32'h3b42332c),
	.w4(32'h3985632c),
	.w5(32'h39560cb4),
	.w6(32'hb7da037f),
	.w7(32'hb95867b5),
	.w8(32'h39cc2d1e),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98c4c63),
	.w1(32'h3b31df74),
	.w2(32'h3ab5c047),
	.w3(32'hbb41c408),
	.w4(32'hbb957c60),
	.w5(32'hbb4ba024),
	.w6(32'hbaa31bae),
	.w7(32'hbb609d0d),
	.w8(32'hbaf457fc),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule