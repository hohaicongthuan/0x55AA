module layer_10_featuremap_176(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb5f9d119),
	.w1(32'h3a40f838),
	.w2(32'h3998b393),
	.w3(32'h38fbf5b8),
	.w4(32'h3a616bd1),
	.w5(32'h3aa577bb),
	.w6(32'h3a8c3944),
	.w7(32'h3a951729),
	.w8(32'h3a887b07),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b755359),
	.w1(32'h3ae766f9),
	.w2(32'h3b2b8dc9),
	.w3(32'h3b5f3621),
	.w4(32'h3a38a8cb),
	.w5(32'h3b1b17d3),
	.w6(32'h3aa52e70),
	.w7(32'h39c906e1),
	.w8(32'h3ad31ca3),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3904d362),
	.w1(32'hb8888e33),
	.w2(32'hb8c65724),
	.w3(32'h38e31e23),
	.w4(32'hb9b28d90),
	.w5(32'hb9c42616),
	.w6(32'hb9bd25b2),
	.w7(32'hb9c00084),
	.w8(32'hb999dae4),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93bc15f),
	.w1(32'hba3ab482),
	.w2(32'hbaca6b7f),
	.w3(32'hb99d0575),
	.w4(32'hba48dd84),
	.w5(32'hbaaa4183),
	.w6(32'h39dfbc58),
	.w7(32'h388be5b7),
	.w8(32'hb7cdb1d2),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba79e3fe),
	.w1(32'h3a592e30),
	.w2(32'h3988db3b),
	.w3(32'hba9c3f02),
	.w4(32'h3a2445cd),
	.w5(32'h3974d844),
	.w6(32'h3a555147),
	.w7(32'h3a6c0ecf),
	.w8(32'h391e8e16),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391a5be5),
	.w1(32'hb925371f),
	.w2(32'hba42d829),
	.w3(32'hb9668657),
	.w4(32'h393fa13a),
	.w5(32'hb95a1259),
	.w6(32'hb8ddcc3e),
	.w7(32'hb9ea44e6),
	.w8(32'hb912e60a),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2416aa),
	.w1(32'h3a7189ac),
	.w2(32'h39beb58c),
	.w3(32'h39d9d062),
	.w4(32'h3a807cb7),
	.w5(32'h39b3b01a),
	.w6(32'h3ae89e8e),
	.w7(32'h3af851d5),
	.w8(32'h39fc4b62),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1c8129),
	.w1(32'hb9586ab9),
	.w2(32'hbaf09e25),
	.w3(32'h3a7dd5e4),
	.w4(32'hbabb4fda),
	.w5(32'hbb274211),
	.w6(32'hb9e47981),
	.w7(32'hba1a2a65),
	.w8(32'hbab397b0),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba70e4d9),
	.w1(32'h3a219df7),
	.w2(32'h3a159847),
	.w3(32'hb861819e),
	.w4(32'h3a8f803b),
	.w5(32'h3a4e9bd8),
	.w6(32'h3a00ad68),
	.w7(32'h3a8b9bbb),
	.w8(32'h3a254bc5),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b26d166),
	.w1(32'h3be9c02c),
	.w2(32'h3c1198d0),
	.w3(32'hba5f228c),
	.w4(32'h3b7687a6),
	.w5(32'h3bed1729),
	.w6(32'hb97f0623),
	.w7(32'h3b309eaa),
	.w8(32'h3be0fcd4),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5371c8),
	.w1(32'h330d6586),
	.w2(32'h39f5d3a0),
	.w3(32'h3a91a7a3),
	.w4(32'hba09e28a),
	.w5(32'hba4be4ac),
	.w6(32'hba5f2000),
	.w7(32'hba849942),
	.w8(32'hba4c4848),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb460019),
	.w1(32'hbb63a8b2),
	.w2(32'hbac03b40),
	.w3(32'hbaf5327a),
	.w4(32'hbacf3916),
	.w5(32'hbaa1a1f2),
	.w6(32'h38f2aa21),
	.w7(32'hba3138b1),
	.w8(32'hba07ff85),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d95d98),
	.w1(32'h3b5284fb),
	.w2(32'h3bba3a33),
	.w3(32'hbb087e19),
	.w4(32'h3adb3e69),
	.w5(32'h3b9e384c),
	.w6(32'hbb270ee9),
	.w7(32'h39f52d1b),
	.w8(32'h3b744456),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h381b38a0),
	.w1(32'hba8278ec),
	.w2(32'hb8993b29),
	.w3(32'hb8b4e13c),
	.w4(32'hb906497e),
	.w5(32'h39d1994b),
	.w6(32'hba675041),
	.w7(32'hbb232145),
	.w8(32'hb9ee9ea0),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38493dba),
	.w1(32'h3b379592),
	.w2(32'h3b8759a9),
	.w3(32'hba985be6),
	.w4(32'h3a83302e),
	.w5(32'h3b44a39d),
	.w6(32'h3a8f418b),
	.w7(32'h3ab0d97a),
	.w8(32'h3b7b22aa),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7d4de0),
	.w1(32'h3b8c0fbb),
	.w2(32'h3bb984e1),
	.w3(32'h3a04e367),
	.w4(32'h3ae398d6),
	.w5(32'h3b8b6b5d),
	.w6(32'hbaa5b157),
	.w7(32'h3a066e85),
	.w8(32'h3b887749),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a7e018),
	.w1(32'hb996d2eb),
	.w2(32'hba4bc3bb),
	.w3(32'h396a79e7),
	.w4(32'hb7dac695),
	.w5(32'hba284be4),
	.w6(32'hba3fad60),
	.w7(32'hba6d5a2f),
	.w8(32'hba4e6b7b),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbdbd68),
	.w1(32'h3a5f9ecf),
	.w2(32'h3a5482a8),
	.w3(32'hbb579bde),
	.w4(32'h399b7c8d),
	.w5(32'hba1e4a5e),
	.w6(32'hba663c7d),
	.w7(32'hb95c7639),
	.w8(32'hbace97cd),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7d7552),
	.w1(32'h39f36741),
	.w2(32'h398019d9),
	.w3(32'hb99fb1d4),
	.w4(32'hb831ff06),
	.w5(32'hb9a45a09),
	.w6(32'hb9da21b5),
	.w7(32'hb94aaef2),
	.w8(32'hba5d4c93),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb91a382e),
	.w1(32'hb9a96d82),
	.w2(32'hb9db3f05),
	.w3(32'hb86c26aa),
	.w4(32'hb96dbde2),
	.w5(32'hb9acdb72),
	.w6(32'hb9a15d7f),
	.w7(32'hb9b6f7e8),
	.w8(32'hb9b1ba1a),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99a9313),
	.w1(32'hb9c49c2c),
	.w2(32'hba6ac2cf),
	.w3(32'hb978a1f4),
	.w4(32'hb8b0d391),
	.w5(32'hba002ae4),
	.w6(32'hb90cd566),
	.w7(32'hb9c30f61),
	.w8(32'hb9fdfdfc),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba88fc6d),
	.w1(32'hbacc57f5),
	.w2(32'hb9fbca22),
	.w3(32'hba2ff0b9),
	.w4(32'hbb0485c4),
	.w5(32'hbae2e11b),
	.w6(32'h3a0d27e4),
	.w7(32'hb93edc04),
	.w8(32'hb89b0787),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb193bff),
	.w1(32'h3b8fc309),
	.w2(32'h3c188bfc),
	.w3(32'hbb71dc57),
	.w4(32'h3aa9622a),
	.w5(32'h3b943c6d),
	.w6(32'hbb70faf3),
	.w7(32'hbb58ba14),
	.w8(32'hb9be51ef),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b80d372),
	.w1(32'h3baab08c),
	.w2(32'h3be921a7),
	.w3(32'h3a421cbf),
	.w4(32'h3b1245d4),
	.w5(32'h3baeb4b2),
	.w6(32'hba95720c),
	.w7(32'h3a7023fe),
	.w8(32'h3bb009a7),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8d552d),
	.w1(32'h3b87420e),
	.w2(32'h3bed9df2),
	.w3(32'h38c1e9f9),
	.w4(32'h3a2bf42d),
	.w5(32'h3b93dd96),
	.w6(32'hbab23808),
	.w7(32'hba72643c),
	.w8(32'h3b90dbdd),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a309ae1),
	.w1(32'h395f7a59),
	.w2(32'h3982753d),
	.w3(32'h39a30a79),
	.w4(32'h3864560c),
	.w5(32'h39429ad9),
	.w6(32'hba1e37ee),
	.w7(32'h382840d3),
	.w8(32'h39f72c61),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3305da),
	.w1(32'hba006621),
	.w2(32'hba247aa1),
	.w3(32'hba5fd6aa),
	.w4(32'hb9c0c68c),
	.w5(32'hba2164c2),
	.w6(32'hb9781a12),
	.w7(32'hb9b86d17),
	.w8(32'hb9e2fad8),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba77065c),
	.w1(32'hbb3366a6),
	.w2(32'hba152e9e),
	.w3(32'hbad994ca),
	.w4(32'hbb014f6d),
	.w5(32'hb9abb0be),
	.w6(32'hbb0ae0b5),
	.w7(32'hbafeeef9),
	.w8(32'h37d74fca),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba77bbcd),
	.w1(32'hbb2efac2),
	.w2(32'hbb0dfdda),
	.w3(32'hba6355b1),
	.w4(32'hbb03ee5a),
	.w5(32'hbb06735a),
	.w6(32'hb9915bd1),
	.w7(32'hbae2cc28),
	.w8(32'hbac16e20),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7b4b07),
	.w1(32'h3b9d37e4),
	.w2(32'h3bccb56c),
	.w3(32'hb9e2a8e3),
	.w4(32'h3abdc4b2),
	.w5(32'h3b9b4347),
	.w6(32'hbb06ba42),
	.w7(32'h39e03223),
	.w8(32'h3b9edd1e),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d4f833),
	.w1(32'hb9b51e5b),
	.w2(32'hba08ba00),
	.w3(32'hb94cf213),
	.w4(32'hb937b6d2),
	.w5(32'hb9c8ac38),
	.w6(32'hb977dfbd),
	.w7(32'hb9c4d942),
	.w8(32'hb9adeb34),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dd6907),
	.w1(32'hb9a08960),
	.w2(32'hb9d9581f),
	.w3(32'hb9cbdf41),
	.w4(32'hb963a7dd),
	.w5(32'hb9c2d4e9),
	.w6(32'hb95f1a88),
	.w7(32'hb9c06015),
	.w8(32'hb9c568ac),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aac6d25),
	.w1(32'h3b12afc8),
	.w2(32'h3b3049f9),
	.w3(32'hb8f67cbb),
	.w4(32'h3a340979),
	.w5(32'h3ad354c6),
	.w6(32'hba86aea5),
	.w7(32'h39a425ba),
	.w8(32'h3ae90e25),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a949bf6),
	.w1(32'h3a44fae7),
	.w2(32'h3aad8ca4),
	.w3(32'h38af0ded),
	.w4(32'h3a21f91b),
	.w5(32'h3ae22803),
	.w6(32'hba859879),
	.w7(32'hb985a04c),
	.w8(32'h3af19cd8),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c26407),
	.w1(32'h3a3c7c9f),
	.w2(32'h38bbdc56),
	.w3(32'hb9324294),
	.w4(32'h3a5ab346),
	.w5(32'h3995f620),
	.w6(32'h39cf53c1),
	.w7(32'h385e019d),
	.w8(32'h394c64c4),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90a4ab8),
	.w1(32'hb920308b),
	.w2(32'hb924cad3),
	.w3(32'h39f92b15),
	.w4(32'h38bbb791),
	.w5(32'hb97678de),
	.w6(32'hb9e695c5),
	.w7(32'h39097402),
	.w8(32'h37d1ff50),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb66f7cb),
	.w1(32'h3a5502c5),
	.w2(32'h3b68af10),
	.w3(32'hbb25e92b),
	.w4(32'h3a11047d),
	.w5(32'h3b0ae381),
	.w6(32'hba5d08e7),
	.w7(32'hba2a85c3),
	.w8(32'hb9ca076c),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b45dfbe),
	.w1(32'hbb8da82e),
	.w2(32'h3bafd3fe),
	.w3(32'hb94220f7),
	.w4(32'hbbadab60),
	.w5(32'h3b4d5585),
	.w6(32'h38d66d20),
	.w7(32'hbb45714c),
	.w8(32'h3b2d03b3),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9cbced),
	.w1(32'hbb0c4ffc),
	.w2(32'h3b29ee11),
	.w3(32'h3b696b47),
	.w4(32'hbb1596e2),
	.w5(32'h3b427c70),
	.w6(32'h3b5045d7),
	.w7(32'hbaea8f42),
	.w8(32'h3b23ea3c),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac4bbd5),
	.w1(32'h3a2a106c),
	.w2(32'h3a32b656),
	.w3(32'h3a068f1a),
	.w4(32'hb90b6f68),
	.w5(32'h39993bcc),
	.w6(32'h3a44df60),
	.w7(32'h39ee3820),
	.w8(32'h39d114f8),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392453bc),
	.w1(32'h392175e2),
	.w2(32'hb8c45875),
	.w3(32'h397d3ecc),
	.w4(32'h393d27ab),
	.w5(32'hb8f16bb1),
	.w6(32'h3986fb72),
	.w7(32'hb8d44611),
	.w8(32'hb9636be3),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9945e68),
	.w1(32'hb9d81c80),
	.w2(32'hb970cf2b),
	.w3(32'hb8c46d4f),
	.w4(32'hb96a6975),
	.w5(32'hb9ff0354),
	.w6(32'hb9845bfc),
	.w7(32'hb9611bc8),
	.w8(32'h33fafe87),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8991af),
	.w1(32'hbac6bcba),
	.w2(32'h3a464852),
	.w3(32'hba9fa6e1),
	.w4(32'hbac72e77),
	.w5(32'h3a44d8b6),
	.w6(32'hba66b4de),
	.w7(32'hbaf61353),
	.w8(32'hb95ca9e4),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b676778),
	.w1(32'h3c1308f0),
	.w2(32'h3bfe50fd),
	.w3(32'h3a093006),
	.w4(32'h3bcdeb6c),
	.w5(32'h3be95bfa),
	.w6(32'h3ab64cea),
	.w7(32'h3b867795),
	.w8(32'h3bd63800),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9522c2),
	.w1(32'h3ba1cffa),
	.w2(32'h3be45ba7),
	.w3(32'h3ab7b1a7),
	.w4(32'h3acd679e),
	.w5(32'h3bad70c0),
	.w6(32'hbaa8a8a9),
	.w7(32'h3a816f66),
	.w8(32'h3bb5d0de),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8f723f),
	.w1(32'h3bd3f2c7),
	.w2(32'h3c0f490f),
	.w3(32'h3863faa5),
	.w4(32'h3b1811a8),
	.w5(32'h3bc76536),
	.w6(32'hba9b532f),
	.w7(32'h3ad812a3),
	.w8(32'h3bd2e87f),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af7cd20),
	.w1(32'h3b43c8c0),
	.w2(32'h3bcd8b06),
	.w3(32'hba23414a),
	.w4(32'hba4f4b41),
	.w5(32'h3b3ee5db),
	.w6(32'hba3d9a43),
	.w7(32'h39e14733),
	.w8(32'h3b7f4665),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a57c0),
	.w1(32'h3a99fd76),
	.w2(32'h3a740e97),
	.w3(32'hbb596918),
	.w4(32'hba1dd9df),
	.w5(32'hbad70884),
	.w6(32'hbb94d560),
	.w7(32'hbb52a476),
	.w8(32'hbb5c2156),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394af329),
	.w1(32'hb91327ee),
	.w2(32'hb91f1fdc),
	.w3(32'hb9a17004),
	.w4(32'hb95df428),
	.w5(32'hb99a3354),
	.w6(32'hb9db892f),
	.w7(32'hb942fc1b),
	.w8(32'hb99b717a),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c586d5),
	.w1(32'h39aa9af5),
	.w2(32'hb991ee6a),
	.w3(32'h3a2af9c4),
	.w4(32'h3a0bf789),
	.w5(32'hb9023bc2),
	.w6(32'h39d54b79),
	.w7(32'h39c705bd),
	.w8(32'h39209d05),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba09565d),
	.w1(32'h3a4a414f),
	.w2(32'h3a1171c7),
	.w3(32'hb99f3b27),
	.w4(32'h3a2b2cc9),
	.w5(32'h39b5f26c),
	.w6(32'h3a43357d),
	.w7(32'h3a197b60),
	.w8(32'h3a32acc6),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38339b37),
	.w1(32'h3b4bab3a),
	.w2(32'h3b8d732d),
	.w3(32'hbac6f687),
	.w4(32'h3a1a0992),
	.w5(32'h3b50988a),
	.w6(32'hbae90281),
	.w7(32'h399fe863),
	.w8(32'h3b21454b),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aadc17c),
	.w1(32'h39bedd17),
	.w2(32'h390206c4),
	.w3(32'h3a4ef25e),
	.w4(32'h39b8a473),
	.w5(32'hb7c9c255),
	.w6(32'h38c0f799),
	.w7(32'hb9c5c932),
	.w8(32'hb95a5b21),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac4b4c4),
	.w1(32'h3b88509f),
	.w2(32'h3b128650),
	.w3(32'hba7bec80),
	.w4(32'h3b6e584a),
	.w5(32'h3b2228fe),
	.w6(32'h3b01a522),
	.w7(32'h3b6b610f),
	.w8(32'h3aa8bff7),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h392cee83),
	.w1(32'hb8e53975),
	.w2(32'hb876f867),
	.w3(32'h39879d66),
	.w4(32'h391c2c53),
	.w5(32'hb8a2776b),
	.w6(32'h3802b2a7),
	.w7(32'hb9f6f952),
	.w8(32'hba2dafc6),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb893858b),
	.w1(32'h392d87e9),
	.w2(32'h3a66584e),
	.w3(32'hb8097e75),
	.w4(32'h3a057cc9),
	.w5(32'h3a770fa6),
	.w6(32'h3843d458),
	.w7(32'h394444ce),
	.w8(32'h3a1e24c6),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1e2459),
	.w1(32'h35083379),
	.w2(32'hb9c78524),
	.w3(32'h3a3072e3),
	.w4(32'h38aae108),
	.w5(32'hb8c5d2b5),
	.w6(32'hb88abfab),
	.w7(32'h38d62d1e),
	.w8(32'h39a94ff2),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397a704a),
	.w1(32'h39e124b0),
	.w2(32'hba01bf13),
	.w3(32'h399a1082),
	.w4(32'h39aa62ae),
	.w5(32'hb90238ef),
	.w6(32'h39d161d2),
	.w7(32'h386d0d28),
	.w8(32'hb8d11a02),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba49104e),
	.w1(32'hba524fc1),
	.w2(32'hb97fc92e),
	.w3(32'hba0db6ba),
	.w4(32'hba17be59),
	.w5(32'h38853c20),
	.w6(32'h3932073c),
	.w7(32'hb9a00933),
	.w8(32'h39b2a8b1),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8556b02),
	.w1(32'hb688c806),
	.w2(32'h392a2e61),
	.w3(32'hb6a25ba7),
	.w4(32'h389eba9e),
	.w5(32'h39045195),
	.w6(32'hb8ba084b),
	.w7(32'hb8ab1aa4),
	.w8(32'hb96aa595),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb168649),
	.w1(32'hb89d9729),
	.w2(32'hb9faf74e),
	.w3(32'hbaae280a),
	.w4(32'h3a2032d0),
	.w5(32'hba0d4506),
	.w6(32'hba97e6f1),
	.w7(32'hb995060c),
	.w8(32'hb8cadfde),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b9d21b),
	.w1(32'h3ac8e18b),
	.w2(32'h3a5568e4),
	.w3(32'h38149338),
	.w4(32'h3a40560e),
	.w5(32'hb898b700),
	.w6(32'hba9f44d7),
	.w7(32'hbaac1d37),
	.w8(32'hbaf66156),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99ab579),
	.w1(32'h3836a7ce),
	.w2(32'h38cddf90),
	.w3(32'hb96ef479),
	.w4(32'hb881208c),
	.w5(32'hb8c359cc),
	.w6(32'h3a0ccb1c),
	.w7(32'hb80e0f9b),
	.w8(32'hb9dac835),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cbbbc0),
	.w1(32'h3aa3aa96),
	.w2(32'h3a56c424),
	.w3(32'hb8047aa4),
	.w4(32'h3abf5835),
	.w5(32'h3a8d31e1),
	.w6(32'h3aa869d2),
	.w7(32'h3a8d33bd),
	.w8(32'h3a9cf20e),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9f900e),
	.w1(32'hb94ed8bd),
	.w2(32'hb9ae5ed2),
	.w3(32'h3abe5a4d),
	.w4(32'hb94fa2c5),
	.w5(32'hb98830e0),
	.w6(32'h3740debb),
	.w7(32'hb93257a7),
	.w8(32'hb920cf64),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb870fc75),
	.w1(32'h3928da72),
	.w2(32'hb96579b6),
	.w3(32'h38861e07),
	.w4(32'h398e72c4),
	.w5(32'hb92d82d9),
	.w6(32'h38f0f100),
	.w7(32'hb88d5555),
	.w8(32'h3946e12a),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a94ec65),
	.w1(32'h3ac15071),
	.w2(32'h3a7b911c),
	.w3(32'h3a5c0fd6),
	.w4(32'h3a0d9ef0),
	.w5(32'hb982b8f0),
	.w6(32'h3a547b35),
	.w7(32'h399ed6e9),
	.w8(32'hba06b0be),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b47ebbf),
	.w1(32'h3b235c6f),
	.w2(32'h3ba3cd67),
	.w3(32'hb89de027),
	.w4(32'h39d13082),
	.w5(32'h3b2966d7),
	.w6(32'hbadd497c),
	.w7(32'hba8dffd9),
	.w8(32'h3b5f2df9),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba20d553),
	.w1(32'h3b196f08),
	.w2(32'h3ba0d4e2),
	.w3(32'hbb0e6747),
	.w4(32'hb98fd795),
	.w5(32'h3b09c61a),
	.w6(32'hbaf28f0c),
	.w7(32'hbaf10cbf),
	.w8(32'h3a53d2cb),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc57fb4),
	.w1(32'h3bd48a6f),
	.w2(32'h3c44fde7),
	.w3(32'h3986509f),
	.w4(32'h3af72626),
	.w5(32'h3c04ede7),
	.w6(32'hbb34e202),
	.w7(32'hb988b87b),
	.w8(32'h3bfa9ded),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396e325b),
	.w1(32'h3a05c064),
	.w2(32'h396d707f),
	.w3(32'h371f2e76),
	.w4(32'h39a94a09),
	.w5(32'h39062824),
	.w6(32'h39e61dd4),
	.w7(32'h39e33a14),
	.w8(32'h39a9a747),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d93d8e),
	.w1(32'hb92c231d),
	.w2(32'hb9d2ccc4),
	.w3(32'h39801904),
	.w4(32'hb626ada3),
	.w5(32'hb9761400),
	.w6(32'hb8f02edc),
	.w7(32'hb80ddd23),
	.w8(32'hb8b39673),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b52c1c),
	.w1(32'hb844f3f2),
	.w2(32'hb903d7dd),
	.w3(32'hb9cfe33b),
	.w4(32'h39165464),
	.w5(32'h389a4a5c),
	.w6(32'h37f74be9),
	.w7(32'h37ea41a1),
	.w8(32'hb8d86bec),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0c3867),
	.w1(32'hba218ef4),
	.w2(32'hbaa4675b),
	.w3(32'hb9825cda),
	.w4(32'hba3e03da),
	.w5(32'hbab83179),
	.w6(32'hba6378e8),
	.w7(32'hba285282),
	.w8(32'hbac680a6),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2b91c9),
	.w1(32'hb9e3a575),
	.w2(32'hba165a5e),
	.w3(32'hba288631),
	.w4(32'hb993fdf8),
	.w5(32'hba249b7e),
	.w6(32'hb9940b89),
	.w7(32'hb9d228d2),
	.w8(32'hb9a3bcae),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0d3f4e),
	.w1(32'hba3c0e6d),
	.w2(32'hb81420ae),
	.w3(32'hba89ee3c),
	.w4(32'h3a390532),
	.w5(32'hb9a6d3d4),
	.w6(32'h3972a54d),
	.w7(32'h39e7ffdb),
	.w8(32'hbab47999),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb88044c),
	.w1(32'hbb2fa533),
	.w2(32'h39ec1efa),
	.w3(32'hbbc03c21),
	.w4(32'hb8a19010),
	.w5(32'hba308928),
	.w6(32'hbb841cf9),
	.w7(32'hbb054a4b),
	.w8(32'hbb1b2eef),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aceda8a),
	.w1(32'h3b443ec7),
	.w2(32'h3bbfbc76),
	.w3(32'hbad01930),
	.w4(32'h3a26150f),
	.w5(32'h3b913e27),
	.w6(32'hbb482406),
	.w7(32'hba10e2a0),
	.w8(32'h3b8021e4),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab5008f),
	.w1(32'h3ac89a09),
	.w2(32'h3aad7d17),
	.w3(32'h3a1b0bea),
	.w4(32'h3a8d9b71),
	.w5(32'h3aaebe7d),
	.w6(32'hb9f47695),
	.w7(32'h386ab066),
	.w8(32'h3a4cc6c6),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3394a3),
	.w1(32'h3aba5892),
	.w2(32'h3a61be57),
	.w3(32'h391a2a6b),
	.w4(32'h3a2af0e9),
	.w5(32'h39bf50f2),
	.w6(32'h39244726),
	.w7(32'h39d7b104),
	.w8(32'h3a31fa05),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ea8686),
	.w1(32'h3acb9a22),
	.w2(32'h3af590ac),
	.w3(32'hba7dfd5b),
	.w4(32'h3988a77e),
	.w5(32'h3ac96c03),
	.w6(32'hba9798e3),
	.w7(32'hb9e01a17),
	.w8(32'h3ad42623),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb02d4d7),
	.w1(32'h3a28ae33),
	.w2(32'h3a114d83),
	.w3(32'hbb150f47),
	.w4(32'h3a097793),
	.w5(32'h3a182457),
	.w6(32'hbac5d793),
	.w7(32'h39a7f814),
	.w8(32'h3a031f48),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94a2345),
	.w1(32'hb964689f),
	.w2(32'hb910dd4c),
	.w3(32'hb8ae6962),
	.w4(32'hb98afc46),
	.w5(32'hb9a0c979),
	.w6(32'hba053df0),
	.w7(32'hba0c4e72),
	.w8(32'hba0690f1),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38707b88),
	.w1(32'hb81cb7c1),
	.w2(32'hb9811ac1),
	.w3(32'hb9811fbf),
	.w4(32'hb7f21add),
	.w5(32'hb961c021),
	.w6(32'h37dc134f),
	.w7(32'h358753ba),
	.w8(32'h38e8c31f),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0ab0e6),
	.w1(32'h3a32bc26),
	.w2(32'h39391063),
	.w3(32'h39c3ff2b),
	.w4(32'hba3b18db),
	.w5(32'hba47b4ba),
	.w6(32'hba1eeaa4),
	.w7(32'hbaa45788),
	.w8(32'hba993c1e),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39291756),
	.w1(32'hb9c90f5a),
	.w2(32'hb9a24490),
	.w3(32'hb9e5adc2),
	.w4(32'hb933966d),
	.w5(32'hb8e96fce),
	.w6(32'hb9b57861),
	.w7(32'hb956ffbb),
	.w8(32'h379ca78a),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b93098f),
	.w1(32'h3b091e21),
	.w2(32'h3b87ca20),
	.w3(32'h3b4a324b),
	.w4(32'h3b087584),
	.w5(32'h3b569329),
	.w6(32'h3a004b23),
	.w7(32'h3a756046),
	.w8(32'h3add0aac),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba446266),
	.w1(32'hbab0070f),
	.w2(32'hba24ca61),
	.w3(32'hb9981683),
	.w4(32'hba4d4bbc),
	.w5(32'hb922fafb),
	.w6(32'hba00db3a),
	.w7(32'hba629348),
	.w8(32'hb9bf4273),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b007bbe),
	.w1(32'h3b84ebc1),
	.w2(32'h3b422e6e),
	.w3(32'h3ab04ffe),
	.w4(32'h3b5576de),
	.w5(32'h3b1c38f1),
	.w6(32'h3b1b3eb5),
	.w7(32'h3b1c1b73),
	.w8(32'h3b4ad601),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h389464ed),
	.w1(32'h3b4a4587),
	.w2(32'h3b1a47c0),
	.w3(32'hb8bc20b0),
	.w4(32'h3b745a28),
	.w5(32'h398f7ea5),
	.w6(32'hb928ede8),
	.w7(32'hb95f545b),
	.w8(32'hbb081939),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba57d30e),
	.w1(32'hbb39749e),
	.w2(32'h3903b3e1),
	.w3(32'hbacd95cb),
	.w4(32'hbb1c2c32),
	.w5(32'hb969d08d),
	.w6(32'hba486a35),
	.w7(32'hbb05349e),
	.w8(32'hba66c2bf),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb00e5a3),
	.w1(32'h3a882724),
	.w2(32'h3b9b2d57),
	.w3(32'hbab38e46),
	.w4(32'h3b0d6f41),
	.w5(32'h3b8169ea),
	.w6(32'h3a0e4a1c),
	.w7(32'h3ae85109),
	.w8(32'h3b8716b9),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8ed767),
	.w1(32'h3940b206),
	.w2(32'h3a88077e),
	.w3(32'h3994f939),
	.w4(32'hb9b3b6d8),
	.w5(32'h3a4fe341),
	.w6(32'hbab3eee2),
	.w7(32'hba61aef2),
	.w8(32'h3a37f135),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b85beeb),
	.w1(32'h3b91f529),
	.w2(32'h3b7117c2),
	.w3(32'h3ad4d679),
	.w4(32'h3a9ef35e),
	.w5(32'h3ab298f4),
	.w6(32'h3a7608f0),
	.w7(32'h3a4e3f19),
	.w8(32'h3b03b411),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0369f1),
	.w1(32'h3b4e532c),
	.w2(32'h3b5d9285),
	.w3(32'h3ae62216),
	.w4(32'h3b4686e9),
	.w5(32'h3b3c7e09),
	.w6(32'h3a8cc64e),
	.w7(32'h3b11322d),
	.w8(32'h3b4aa97d),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b04737a),
	.w1(32'h3b220b4f),
	.w2(32'h3b916109),
	.w3(32'hba9d21f7),
	.w4(32'h3a2a4d8d),
	.w5(32'h3b3ed222),
	.w6(32'hb8e0dba7),
	.w7(32'h3af053f6),
	.w8(32'h3b45f7e4),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a069908),
	.w1(32'hba8e495b),
	.w2(32'hbab91fbe),
	.w3(32'h3a3fdee8),
	.w4(32'hb9a684e3),
	.w5(32'hba425cad),
	.w6(32'hb9f6f73d),
	.w7(32'hba3906bb),
	.w8(32'hba4fde4b),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39da0ad6),
	.w1(32'h3b8c869b),
	.w2(32'h3bb665fe),
	.w3(32'hba2382db),
	.w4(32'h3abc978f),
	.w5(32'h3b60a9ca),
	.w6(32'hba80d3cc),
	.w7(32'h391694a4),
	.w8(32'h3b24a8e9),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba28e53a),
	.w1(32'h3abf9f0d),
	.w2(32'h3b774344),
	.w3(32'h3989ae31),
	.w4(32'h3afe4e91),
	.w5(32'h3b650f3c),
	.w6(32'h3a2b4363),
	.w7(32'h3ad8c597),
	.w8(32'h3b246be3),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9c21bd),
	.w1(32'hbadc37f7),
	.w2(32'hbae63b88),
	.w3(32'hbb68658f),
	.w4(32'h3b0d722b),
	.w5(32'hb6d9705f),
	.w6(32'hbace773b),
	.w7(32'hb99b1d5e),
	.w8(32'hbb106cee),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcc9b9c),
	.w1(32'h3a93a561),
	.w2(32'h3c1d1c0f),
	.w3(32'h3bf81d1d),
	.w4(32'h3b11023d),
	.w5(32'h3bf0daf6),
	.w6(32'h3b869af0),
	.w7(32'h3a0ba0ff),
	.w8(32'h3baa14fd),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bad6ee9),
	.w1(32'h3c0149b9),
	.w2(32'h3c188980),
	.w3(32'h3a270fa5),
	.w4(32'h3b9c4640),
	.w5(32'h3bf43394),
	.w6(32'h39ac5e29),
	.w7(32'h3b5b0bb3),
	.w8(32'h3c081dd5),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8b08e35),
	.w1(32'h3aa1d5f4),
	.w2(32'h3afab35f),
	.w3(32'hb82ad911),
	.w4(32'h3aa00a73),
	.w5(32'h3945fce0),
	.w6(32'h3a3c6eb8),
	.w7(32'hb997837c),
	.w8(32'hbaaa94e8),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba511b48),
	.w1(32'h3907cc36),
	.w2(32'hb93c9b9e),
	.w3(32'h3696adc5),
	.w4(32'h39d14a90),
	.w5(32'hb8c8a00e),
	.w6(32'h384a1af0),
	.w7(32'h3861dfd3),
	.w8(32'hb965871a),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba5f731),
	.w1(32'hbb186970),
	.w2(32'hb98960fd),
	.w3(32'hbba3533a),
	.w4(32'hb9fd7a39),
	.w5(32'hb8802ac6),
	.w6(32'hbaa533fd),
	.w7(32'h39721a4c),
	.w8(32'hbb7687b2),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99c815e),
	.w1(32'hbadf502a),
	.w2(32'h3b16b9c0),
	.w3(32'hbb29b318),
	.w4(32'hba9f71ee),
	.w5(32'h3acb15a5),
	.w6(32'hbb7293b9),
	.w7(32'hba0fe520),
	.w8(32'h3a83b868),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d87436),
	.w1(32'hb99102f5),
	.w2(32'hb8ac7253),
	.w3(32'hb9bfae5f),
	.w4(32'hba17478d),
	.w5(32'hba23375f),
	.w6(32'hba00233a),
	.w7(32'hba09e9e9),
	.w8(32'hba075a7b),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4e71ea),
	.w1(32'h3a021f23),
	.w2(32'h39dac1bc),
	.w3(32'h38af7f02),
	.w4(32'h3930140f),
	.w5(32'h39d69736),
	.w6(32'h3980e75a),
	.w7(32'hb9ab7b9a),
	.w8(32'hb94cc638),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1e7d0e),
	.w1(32'h3b955a37),
	.w2(32'h3baac809),
	.w3(32'hba89b6f4),
	.w4(32'h3abfd5f0),
	.w5(32'h3b8084e6),
	.w6(32'hbae66845),
	.w7(32'h390b74ad),
	.w8(32'h3b5fa6e5),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b55aaaa),
	.w1(32'h3bb35aaf),
	.w2(32'h3bd3af93),
	.w3(32'hb818e273),
	.w4(32'h3b1a6fab),
	.w5(32'h3bab79ff),
	.w6(32'hba7309c4),
	.w7(32'h3ae3af06),
	.w8(32'h3ba6688b),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b59bc19),
	.w1(32'h3b015a2f),
	.w2(32'h3b29630b),
	.w3(32'h3af2dfbb),
	.w4(32'hb8757b27),
	.w5(32'h3a7a7772),
	.w6(32'h396942bd),
	.w7(32'hb9a75589),
	.w8(32'h392708fb),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b015c0a),
	.w1(32'h3b25d9e0),
	.w2(32'h3b79e638),
	.w3(32'h3a96ff33),
	.w4(32'h3a70abe9),
	.w5(32'h3b51650a),
	.w6(32'hb965f848),
	.w7(32'h3a770a5f),
	.w8(32'h3b0b0ed2),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba442a50),
	.w1(32'hba82fd90),
	.w2(32'h3a492be6),
	.w3(32'hba3e4807),
	.w4(32'hba47398f),
	.w5(32'h39f95e3c),
	.w6(32'hb9f2ebf4),
	.w7(32'hba873e8d),
	.w8(32'h3a1bc175),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c3b0f6),
	.w1(32'h3a9b33e4),
	.w2(32'h3b022b9f),
	.w3(32'hb9e8d24d),
	.w4(32'h3ad2adfc),
	.w5(32'h3af6ead0),
	.w6(32'hbac2e958),
	.w7(32'h3919fd86),
	.w8(32'h3a842c96),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1e146a),
	.w1(32'h3b38de96),
	.w2(32'h3b7b94e2),
	.w3(32'h3911181d),
	.w4(32'h3a15f1a6),
	.w5(32'h3b374aea),
	.w6(32'hba977747),
	.w7(32'h399ba0bf),
	.w8(32'h3b229cd9),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3709ba),
	.w1(32'hba2911b5),
	.w2(32'hba92ae1b),
	.w3(32'hba202524),
	.w4(32'hb8aa20d5),
	.w5(32'hba1524d2),
	.w6(32'hb9b30549),
	.w7(32'hba68afae),
	.w8(32'hba2b45c4),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5949f8),
	.w1(32'hb9b74552),
	.w2(32'hba182d35),
	.w3(32'hb99a253e),
	.w4(32'hb902e1f4),
	.w5(32'hb9a08544),
	.w6(32'hb9cdbabc),
	.w7(32'hba29715a),
	.w8(32'hba0604e6),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e9625a),
	.w1(32'hb9fb77d2),
	.w2(32'hba4ffb43),
	.w3(32'hb933f744),
	.w4(32'hb8dac393),
	.w5(32'hb9f49b77),
	.w6(32'hb9c58686),
	.w7(32'hba4ceb00),
	.w8(32'hba2115e0),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba14d5dd),
	.w1(32'h3a1a0976),
	.w2(32'h38dc45c6),
	.w3(32'hb962b5d6),
	.w4(32'hb92ed314),
	.w5(32'hba102881),
	.w6(32'h39eed953),
	.w7(32'h3892575a),
	.w8(32'hb6d97b9a),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b33bc2d),
	.w1(32'h3b5e2ff1),
	.w2(32'h3b8623cf),
	.w3(32'hb755f8e4),
	.w4(32'h3aa8fde4),
	.w5(32'h3b5d0d5b),
	.w6(32'hba26c6ac),
	.w7(32'h3a30defb),
	.w8(32'h3b4a8be6),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e2b065),
	.w1(32'hba763ea8),
	.w2(32'hba490e4c),
	.w3(32'hba026cf1),
	.w4(32'hba45bafd),
	.w5(32'hba6e9ebd),
	.w6(32'hba4559e5),
	.w7(32'hba8625be),
	.w8(32'hba3b2a07),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0d1329),
	.w1(32'hba248f9d),
	.w2(32'h38c8ac33),
	.w3(32'hbac23ad8),
	.w4(32'hb86ab7f4),
	.w5(32'hba0104de),
	.w6(32'hb9ae854b),
	.w7(32'h392dd6e7),
	.w8(32'hb9e93102),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b341d75),
	.w1(32'h3b2de3a6),
	.w2(32'h3ba3cbb1),
	.w3(32'hb9933290),
	.w4(32'h3a9e6d36),
	.w5(32'h3bc918ba),
	.w6(32'hba7aac21),
	.w7(32'h3a958de2),
	.w8(32'h3b97a304),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a141ab),
	.w1(32'h3aad3773),
	.w2(32'h3a8839cc),
	.w3(32'hb98d9fdc),
	.w4(32'h3a748f14),
	.w5(32'h3a4f2331),
	.w6(32'h3ad4d9a5),
	.w7(32'h3b0736a0),
	.w8(32'h3ab58618),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1c9b8a),
	.w1(32'hb89f9836),
	.w2(32'hba439bad),
	.w3(32'h3aa5c57a),
	.w4(32'h38ddcfca),
	.w5(32'hb9d562b8),
	.w6(32'h39d164ff),
	.w7(32'hb8fd5e1f),
	.w8(32'hb93da5df),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92bf94f),
	.w1(32'hba0d7091),
	.w2(32'hba514114),
	.w3(32'h35ce9f73),
	.w4(32'hb9b59cbc),
	.w5(32'hba24f5f7),
	.w6(32'hba080521),
	.w7(32'hba3053f0),
	.w8(32'hba0c040b),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c0a10c),
	.w1(32'h3b7806e7),
	.w2(32'h3b35d5c9),
	.w3(32'h399ec45f),
	.w4(32'h3a51db72),
	.w5(32'h39df7ec1),
	.w6(32'h39f5c317),
	.w7(32'h39b7d2fa),
	.w8(32'hbb8efbbe),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3db13a),
	.w1(32'h3b0e162f),
	.w2(32'h3b9fa01d),
	.w3(32'hbb86fa83),
	.w4(32'h3a35e589),
	.w5(32'h3b6fc67b),
	.w6(32'hbb29290d),
	.w7(32'h3b11ae82),
	.w8(32'h3aaccdfc),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9584af),
	.w1(32'hbb5d3cda),
	.w2(32'h3ba5d7bc),
	.w3(32'h3b22ef96),
	.w4(32'hbbe291af),
	.w5(32'h3a448ad0),
	.w6(32'hbabe8089),
	.w7(32'h3c1f5524),
	.w8(32'h3beb6acc),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b86a2d0),
	.w1(32'hbaef51de),
	.w2(32'hbb277b85),
	.w3(32'hba9b85f8),
	.w4(32'hbadd55e3),
	.w5(32'hbb1e6b5b),
	.w6(32'hbac93615),
	.w7(32'hbb1c73fa),
	.w8(32'hbafa45cb),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac52987),
	.w1(32'hbae28b6c),
	.w2(32'hbada141b),
	.w3(32'hbad2899f),
	.w4(32'hbabde6e9),
	.w5(32'hbb05f302),
	.w6(32'hbad0601e),
	.w7(32'hbb32d702),
	.w8(32'hb9fa4d11),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf247ab),
	.w1(32'h3b1463d4),
	.w2(32'hba4fc379),
	.w3(32'hbaa10177),
	.w4(32'h3a1fac0c),
	.w5(32'h383a54f8),
	.w6(32'hbb6b809c),
	.w7(32'hbbc3c7cb),
	.w8(32'hbb2f3d19),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5cb929),
	.w1(32'h3b9523e6),
	.w2(32'h3baa8b0e),
	.w3(32'h386a1d9d),
	.w4(32'h3b3aeb3d),
	.w5(32'h3bba25f4),
	.w6(32'hb89e321a),
	.w7(32'h3a06ae6b),
	.w8(32'hba8bc3db),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b196907),
	.w1(32'h3bffe1a7),
	.w2(32'h3c12532c),
	.w3(32'h3b8e1f98),
	.w4(32'h3baea88f),
	.w5(32'h3c0f1b21),
	.w6(32'h3b4a170a),
	.w7(32'h3bee1406),
	.w8(32'h3c1286ba),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baf0fda),
	.w1(32'hbb8aeb81),
	.w2(32'hbb5ad70d),
	.w3(32'h3ba7c30d),
	.w4(32'hbb32feb1),
	.w5(32'hbb394948),
	.w6(32'hbb947526),
	.w7(32'hbb86702c),
	.w8(32'hbb3c9d3b),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab0fe26),
	.w1(32'h3b37fca7),
	.w2(32'h3be757ad),
	.w3(32'hbb3c129c),
	.w4(32'hba902277),
	.w5(32'h3ba9d58a),
	.w6(32'hbb6159d5),
	.w7(32'h39f0c329),
	.w8(32'h3ad06c88),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b39817c),
	.w1(32'h3b075673),
	.w2(32'h3beae71b),
	.w3(32'h3a814727),
	.w4(32'h3aaf5d8d),
	.w5(32'h3bf0fbd6),
	.w6(32'hbaced98b),
	.w7(32'h3b6a73d3),
	.w8(32'hb975c646),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5aa768),
	.w1(32'hbbb4bd28),
	.w2(32'hbbbd1000),
	.w3(32'h3a64497c),
	.w4(32'hbb783c97),
	.w5(32'hbbaa1c9c),
	.w6(32'hbbe4528e),
	.w7(32'hbc0ae276),
	.w8(32'hbb9e44ef),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf1b3cb),
	.w1(32'h3ba35562),
	.w2(32'h3be8f6ff),
	.w3(32'hbb014d8f),
	.w4(32'hbba1a3db),
	.w5(32'hbba38271),
	.w6(32'h3b92a92c),
	.w7(32'h3b89fd5b),
	.w8(32'h3c041626),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf70481),
	.w1(32'h3a2e2b61),
	.w2(32'h3b8dd978),
	.w3(32'hbbcbbdb7),
	.w4(32'h3a51888f),
	.w5(32'h3bb1659a),
	.w6(32'hbc15fde8),
	.w7(32'hbbcef4a3),
	.w8(32'hbb090bb3),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeca001),
	.w1(32'h3b27bd56),
	.w2(32'h3b409831),
	.w3(32'h3b55f67c),
	.w4(32'hba560c90),
	.w5(32'h3906bdba),
	.w6(32'h3a914617),
	.w7(32'h3b364ff2),
	.w8(32'h39f20703),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd34e18),
	.w1(32'hb8e5e571),
	.w2(32'h3bf6f063),
	.w3(32'hbaca2c81),
	.w4(32'hbb9e3e74),
	.w5(32'h3bc7ece3),
	.w6(32'hbc19de9d),
	.w7(32'hbb22ab1b),
	.w8(32'h39a2b32e),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b109d6d),
	.w1(32'h3c0c86df),
	.w2(32'h3bd2abb0),
	.w3(32'hb9a1270e),
	.w4(32'h3b5e5f5c),
	.w5(32'h3b89fb5c),
	.w6(32'hba9b90df),
	.w7(32'hbb058a40),
	.w8(32'hbb5fa28f),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4366a9),
	.w1(32'h3a292e4d),
	.w2(32'h3b9336b6),
	.w3(32'h3a19f788),
	.w4(32'h3aa5f072),
	.w5(32'h3ba3d1ce),
	.w6(32'hb9c4101f),
	.w7(32'h3b41e3da),
	.w8(32'h3a56eaac),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4641a6),
	.w1(32'h38eb4617),
	.w2(32'hbac46fcf),
	.w3(32'h3b5bab03),
	.w4(32'hbab3b0da),
	.w5(32'hbb6b25a6),
	.w6(32'h390f8627),
	.w7(32'hbb090945),
	.w8(32'hbb39ba27),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf508d3),
	.w1(32'hbc05e6e5),
	.w2(32'hbbe0043a),
	.w3(32'hbb4fcd79),
	.w4(32'hbc0e6533),
	.w5(32'hbbdeed39),
	.w6(32'hbc016a94),
	.w7(32'hbc06f7a5),
	.w8(32'hbbb7ac4c),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5eec84),
	.w1(32'h3b087e8e),
	.w2(32'h3b08a8ff),
	.w3(32'hbbbd2e96),
	.w4(32'h393238e6),
	.w5(32'h3a564724),
	.w6(32'h3ac1daad),
	.w7(32'h3a0f0d42),
	.w8(32'h3aef7a33),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d2a3b9),
	.w1(32'h3aedef12),
	.w2(32'h3bdb5b2f),
	.w3(32'hbabd5069),
	.w4(32'hba0eaf02),
	.w5(32'h3bbb2d0e),
	.w6(32'hbb7b8b00),
	.w7(32'h3a993495),
	.w8(32'h3ae5c8c2),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4b36ca),
	.w1(32'h3ad9a291),
	.w2(32'h3ba3c395),
	.w3(32'hba5862c0),
	.w4(32'hbaf81595),
	.w5(32'h3aa3244b),
	.w6(32'hbb2719f0),
	.w7(32'h3a8590ab),
	.w8(32'hbb857ad8),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b722ed0),
	.w1(32'h3b1f8517),
	.w2(32'h3b39a804),
	.w3(32'h3a069d13),
	.w4(32'h3b5d8a6f),
	.w5(32'h3ba969ed),
	.w6(32'hbb425091),
	.w7(32'hba17393d),
	.w8(32'hb9091eb0),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba49b2dd),
	.w1(32'h3ba3a213),
	.w2(32'h3b11891e),
	.w3(32'h3a5986ee),
	.w4(32'h3ba25557),
	.w5(32'h3b5b7973),
	.w6(32'h3b776921),
	.w7(32'h3ad5e225),
	.w8(32'h3bbc9c59),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5e6be3),
	.w1(32'h3a9385fc),
	.w2(32'h3ba69dfc),
	.w3(32'h3b2ce07f),
	.w4(32'hba3af122),
	.w5(32'h3b6290b4),
	.w6(32'hbb6fee39),
	.w7(32'h3af409d2),
	.w8(32'hb8f845bc),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b617ab0),
	.w1(32'h3bed69d9),
	.w2(32'h3c1a9b25),
	.w3(32'hba772d02),
	.w4(32'h3b8b4820),
	.w5(32'h3bacf9ef),
	.w6(32'h3a6e5842),
	.w7(32'h3b8625fc),
	.w8(32'h3bf4247c),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bec2daf),
	.w1(32'hbb569cad),
	.w2(32'hbb80b90d),
	.w3(32'h3b8660e8),
	.w4(32'h3b700aac),
	.w5(32'h3b0d41b7),
	.w6(32'hbbcdd502),
	.w7(32'hbc09dc9d),
	.w8(32'hbbab63fb),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3a3162),
	.w1(32'hbaa1ddd4),
	.w2(32'h39cb90da),
	.w3(32'h3af7514c),
	.w4(32'hbb0ee18e),
	.w5(32'hba5f6305),
	.w6(32'hbb0652b5),
	.w7(32'hba145405),
	.w8(32'hbaaaf953),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398bee34),
	.w1(32'h3b8292eb),
	.w2(32'h3b93b3a2),
	.w3(32'hbb4f621c),
	.w4(32'h3b55952c),
	.w5(32'h3b358b30),
	.w6(32'hbaf90b87),
	.w7(32'hba2b4976),
	.w8(32'h3b12e804),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcb93b4),
	.w1(32'h3bd90b37),
	.w2(32'h3b812569),
	.w3(32'h3b9f08db),
	.w4(32'h3bbf06ca),
	.w5(32'h3b398412),
	.w6(32'h3c250e30),
	.w7(32'h3ba76f59),
	.w8(32'h3a403a2d),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba86fa73),
	.w1(32'hb983adfe),
	.w2(32'hb9ef2c47),
	.w3(32'hbb52346e),
	.w4(32'h39be1551),
	.w5(32'hba613bd5),
	.w6(32'h3a69b013),
	.w7(32'hba7b0d53),
	.w8(32'hbb23f089),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb41eb7a),
	.w1(32'h3a4d5991),
	.w2(32'h3b10e966),
	.w3(32'hbb4bc651),
	.w4(32'hbad16454),
	.w5(32'hbaab8e87),
	.w6(32'hbab81253),
	.w7(32'h39e63cf0),
	.w8(32'hbb3d89ac),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9914ef1),
	.w1(32'hbaf890c9),
	.w2(32'hba927e79),
	.w3(32'hbb2b0822),
	.w4(32'hbb8a9fb5),
	.w5(32'hbb51c328),
	.w6(32'hbb431157),
	.w7(32'hbacaf395),
	.w8(32'hbb3413eb),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2402a7),
	.w1(32'hbb87698a),
	.w2(32'h3b613ad3),
	.w3(32'hbb8f18b6),
	.w4(32'hbb86481f),
	.w5(32'h3a67f01f),
	.w6(32'hbb7fd100),
	.w7(32'h3ad74fe3),
	.w8(32'h3b30e13e),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ab73a6),
	.w1(32'h3a64c2d9),
	.w2(32'hbbc741aa),
	.w3(32'hbb1664f1),
	.w4(32'h3b5eb277),
	.w5(32'hbbc02618),
	.w6(32'h39ebf284),
	.w7(32'hbb87f94f),
	.w8(32'hbbc791f9),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbd66b6),
	.w1(32'h3af1fb86),
	.w2(32'h3b5d5e67),
	.w3(32'hbbca6300),
	.w4(32'h3a1132ab),
	.w5(32'h3b193108),
	.w6(32'hbad4db98),
	.w7(32'hb9a9e1d7),
	.w8(32'h3b43d023),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a891e70),
	.w1(32'h3aa2eafa),
	.w2(32'h3b24d693),
	.w3(32'h3aee43b9),
	.w4(32'hbaa15292),
	.w5(32'hba85d8f2),
	.w6(32'hbad5478e),
	.w7(32'h3a040fca),
	.w8(32'hba5f1c53),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a228c84),
	.w1(32'h3ba8eaea),
	.w2(32'h3b75a8ac),
	.w3(32'hbb159d9d),
	.w4(32'h3b649c6a),
	.w5(32'h3b3198b1),
	.w6(32'h3b9212a3),
	.w7(32'h3b92d503),
	.w8(32'h3bc25227),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc1eaf5),
	.w1(32'hbb9e96d2),
	.w2(32'hbbb5af1c),
	.w3(32'h3b9e715d),
	.w4(32'hbb910957),
	.w5(32'hbba36485),
	.w6(32'hbb85d9a0),
	.w7(32'hbba89521),
	.w8(32'hbb85f09c),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9cf925),
	.w1(32'h399ba1d5),
	.w2(32'h3b45a0c7),
	.w3(32'hbb76305a),
	.w4(32'hbacd3d0a),
	.w5(32'h3aea8507),
	.w6(32'hbb0b03b8),
	.w7(32'h3ab61ad4),
	.w8(32'hb9a652e9),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bca9daf),
	.w1(32'h3b0c3ccc),
	.w2(32'h3ad5517f),
	.w3(32'h3b122512),
	.w4(32'hba72579e),
	.w5(32'h39ba268d),
	.w6(32'h39da8cd3),
	.w7(32'hbad185d7),
	.w8(32'h3a28d9f8),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba446968),
	.w1(32'h3b378c6d),
	.w2(32'h3b338250),
	.w3(32'hb9b659ce),
	.w4(32'h3af1c843),
	.w5(32'h3a1de693),
	.w6(32'hb93eb6c3),
	.w7(32'hba0b9c64),
	.w8(32'h3af28ab5),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb11e053),
	.w1(32'hbb2478a9),
	.w2(32'hba662a99),
	.w3(32'hbab95afc),
	.w4(32'hbb822b8c),
	.w5(32'hbb8b40f5),
	.w6(32'hba935b2d),
	.w7(32'hba87f7fa),
	.w8(32'h370a344c),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b13091e),
	.w1(32'h3a9ed01d),
	.w2(32'h3b96e05b),
	.w3(32'hbb88c313),
	.w4(32'hbb4d7a29),
	.w5(32'h3af477b7),
	.w6(32'hbb4b1c1b),
	.w7(32'h3a20e3a9),
	.w8(32'h3b8c0b2e),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6c92f9),
	.w1(32'hbc09416e),
	.w2(32'hbbbd820c),
	.w3(32'hbb0248ca),
	.w4(32'hbbc683aa),
	.w5(32'hbb98a5f7),
	.w6(32'hbc27755d),
	.w7(32'hbc2ebb01),
	.w8(32'hbb6c0be5),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6703bc),
	.w1(32'hbc4c1752),
	.w2(32'hbc20d4cc),
	.w3(32'hb8d34228),
	.w4(32'hbc3c95af),
	.w5(32'hbc1e3a11),
	.w6(32'hbc4acba4),
	.w7(32'hbc5330d6),
	.w8(32'hbc2fe761),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc428aaf),
	.w1(32'hbbbd96f3),
	.w2(32'hbb988d15),
	.w3(32'hbc41912e),
	.w4(32'hbbcb139e),
	.w5(32'hbbb4fa89),
	.w6(32'hbbddacb9),
	.w7(32'hbbfe9c9c),
	.w8(32'hbba4888f),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb7698c),
	.w1(32'h3b07942f),
	.w2(32'h3b8d0096),
	.w3(32'hbbb9e4c9),
	.w4(32'h3abc868a),
	.w5(32'h3bba0686),
	.w6(32'hbbd5346c),
	.w7(32'hbb555c3f),
	.w8(32'hb9bbfb3c),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ea7195),
	.w1(32'h3bcb2da4),
	.w2(32'h3b8a25e8),
	.w3(32'h3acc9094),
	.w4(32'h3b8ad211),
	.w5(32'h3aa11c0e),
	.w6(32'h3bdcdff8),
	.w7(32'h3b9aec61),
	.w8(32'hb8e80bea),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8e21ba5),
	.w1(32'hba1b3029),
	.w2(32'hbaab70c4),
	.w3(32'hbb3b851c),
	.w4(32'hbb06084d),
	.w5(32'hbb1d2fa1),
	.w6(32'hba8e782b),
	.w7(32'h3797dfaa),
	.w8(32'hba7f305c),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6005f5),
	.w1(32'hb9ff6bf4),
	.w2(32'h3b2ab080),
	.w3(32'hbb13beb6),
	.w4(32'hbb06b4d2),
	.w5(32'h3ad6bac4),
	.w6(32'hbb584521),
	.w7(32'h37e79286),
	.w8(32'hba87fef0),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b26e812),
	.w1(32'hbc2a260a),
	.w2(32'hbc347dd1),
	.w3(32'h3a2aba31),
	.w4(32'hbc2725e0),
	.w5(32'hbc2c744e),
	.w6(32'hbc306598),
	.w7(32'hbc4836bf),
	.w8(32'hbc201a3c),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2fe0f8),
	.w1(32'hbc04c201),
	.w2(32'h3bd0c3d5),
	.w3(32'hbc1f7770),
	.w4(32'hbbc7b30a),
	.w5(32'h3b8dc2c8),
	.w6(32'hbc4689ec),
	.w7(32'hb9b124af),
	.w8(32'hbaa8c6d0),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd8892f),
	.w1(32'h3bcdf616),
	.w2(32'h3c186d7d),
	.w3(32'h3b34ea68),
	.w4(32'h3ba325f0),
	.w5(32'h3c022dcb),
	.w6(32'h3b678e90),
	.w7(32'h3bf3ef10),
	.w8(32'h3c1b82df),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1d5914),
	.w1(32'h3b3e722a),
	.w2(32'hb9d2393f),
	.w3(32'h3c099d5f),
	.w4(32'h3b1a0fcf),
	.w5(32'h3976cdf8),
	.w6(32'h3ac942cf),
	.w7(32'hb98c717d),
	.w8(32'h3a9721f2),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d1f31d),
	.w1(32'h3b4ef655),
	.w2(32'h3ac4cca8),
	.w3(32'h3b14aac9),
	.w4(32'h3b6dd269),
	.w5(32'h3b1744a3),
	.w6(32'h3b6c8cef),
	.w7(32'h3b32fab1),
	.w8(32'h3ba27f0c),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8072b4),
	.w1(32'h3b001c6e),
	.w2(32'h3a1854ef),
	.w3(32'h3b9754a2),
	.w4(32'h3aa3411f),
	.w5(32'hbaf153f8),
	.w6(32'h399e430d),
	.w7(32'hbb07d913),
	.w8(32'h39e8c0dd),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a375022),
	.w1(32'hbbd5e303),
	.w2(32'hbbb68328),
	.w3(32'hba0c1c70),
	.w4(32'hbbd652fe),
	.w5(32'hbbbdba4a),
	.w6(32'hbbe3a1fd),
	.w7(32'hbc1a1fde),
	.w8(32'hbbda2388),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc23f216),
	.w1(32'h3c0199ec),
	.w2(32'h3ab340e3),
	.w3(32'hbc16d481),
	.w4(32'h3bdfa0d4),
	.w5(32'h3b08f8b0),
	.w6(32'h3b9d9572),
	.w7(32'hba4b3802),
	.w8(32'hb9c7dea8),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9cbff6),
	.w1(32'hbb5a129b),
	.w2(32'hbb977c21),
	.w3(32'hba658206),
	.w4(32'hbb3f1c52),
	.w5(32'hbb76d324),
	.w6(32'hbb718c99),
	.w7(32'hbb9aac5d),
	.w8(32'hbb78da2e),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc24b84a),
	.w1(32'h3b0c70d5),
	.w2(32'h3bb440ce),
	.w3(32'hbc116c4c),
	.w4(32'h3abc6a17),
	.w5(32'h3b9f1c98),
	.w6(32'hbbf1e01d),
	.w7(32'h3af40eae),
	.w8(32'h3b2babe9),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c15f244),
	.w1(32'h3b97fe21),
	.w2(32'h3b96c24b),
	.w3(32'h3b80531b),
	.w4(32'h3adf675a),
	.w5(32'h3b3763ad),
	.w6(32'h3b66b281),
	.w7(32'h3a43c77a),
	.w8(32'h3b08b427),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5c5e5e),
	.w1(32'h3889be2e),
	.w2(32'h3ba3162c),
	.w3(32'hb9130e40),
	.w4(32'hbb58e106),
	.w5(32'h3a91b05b),
	.w6(32'hb75ad374),
	.w7(32'h3b7961b0),
	.w8(32'h3a976822),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b65cbee),
	.w1(32'h3ad2fcd2),
	.w2(32'h3c08c8e3),
	.w3(32'h39594ae0),
	.w4(32'h3b0e5a53),
	.w5(32'h3c06a00c),
	.w6(32'h3ba68bc7),
	.w7(32'h3c211fd1),
	.w8(32'hba309c7f),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb50198e),
	.w1(32'hbbc94033),
	.w2(32'hbba5a2be),
	.w3(32'hbb896002),
	.w4(32'hbb91aee6),
	.w5(32'hbb879297),
	.w6(32'hbbe195f9),
	.w7(32'hbbf8af60),
	.w8(32'hbb43f111),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb015043),
	.w1(32'h38ac439d),
	.w2(32'h390c7769),
	.w3(32'h39348c21),
	.w4(32'hb967d7e8),
	.w5(32'h386b11b4),
	.w6(32'h3a85c341),
	.w7(32'h3a5c6dac),
	.w8(32'h3b1d164b),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af813a7),
	.w1(32'h3b6f9836),
	.w2(32'hbab3d685),
	.w3(32'h3ae0f6b4),
	.w4(32'h3b3e300f),
	.w5(32'hbab4f4e3),
	.w6(32'h3b3474df),
	.w7(32'hb98a5160),
	.w8(32'hbb448858),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb36f029),
	.w1(32'h3b874280),
	.w2(32'h3b7739db),
	.w3(32'hbb6a1e17),
	.w4(32'h3b6a804d),
	.w5(32'h3aecde8c),
	.w6(32'h3b3d63a3),
	.w7(32'h3b1cab72),
	.w8(32'hb9dbac4e),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aad670d),
	.w1(32'h3b81074c),
	.w2(32'h3aac2ced),
	.w3(32'hbb285c00),
	.w4(32'h3b1c6055),
	.w5(32'h3a1988d5),
	.w6(32'h3aa08299),
	.w7(32'h3aa306d4),
	.w8(32'h3b7a7642),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadb3c8e),
	.w1(32'h39a9ee09),
	.w2(32'h3ba0a03d),
	.w3(32'hba1c18cc),
	.w4(32'hba729963),
	.w5(32'h3b379326),
	.w6(32'hbac86899),
	.w7(32'h3af05dd3),
	.w8(32'h3b07b357),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8a7301),
	.w1(32'hbc63b55d),
	.w2(32'hbc399da8),
	.w3(32'h3a548f56),
	.w4(32'hbc6886ed),
	.w5(32'hbc4c9d14),
	.w6(32'hbc939d13),
	.w7(32'hbc929473),
	.w8(32'hbc48d747),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc782d0a),
	.w1(32'hbb9cc44e),
	.w2(32'hbb588333),
	.w3(32'hbc85843b),
	.w4(32'hbbabf85a),
	.w5(32'hbb563a11),
	.w6(32'hbba269e7),
	.w7(32'hbb841ba4),
	.w8(32'hbb4a49e8),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c6ea3),
	.w1(32'h3aa89123),
	.w2(32'h3ab8c5fb),
	.w3(32'hbb726e7d),
	.w4(32'hbab86454),
	.w5(32'hb96c26ec),
	.w6(32'hb9ab7d5d),
	.w7(32'h3a92ac71),
	.w8(32'hba996a10),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6e7080),
	.w1(32'hb9f6875c),
	.w2(32'h3b1adf40),
	.w3(32'hbab1908f),
	.w4(32'hbae79c78),
	.w5(32'h3a8a33b8),
	.w6(32'hbb243377),
	.w7(32'h3aa16050),
	.w8(32'hba7ddb7c),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b201085),
	.w1(32'hbaa59497),
	.w2(32'h3a7ffa69),
	.w3(32'h3a5ffd86),
	.w4(32'hbb97e33d),
	.w5(32'hbb5000ed),
	.w6(32'hbb31f556),
	.w7(32'h39f2d0cd),
	.w8(32'hba8f7238),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa1a72b),
	.w1(32'h3ab0d9d7),
	.w2(32'h3b93d9c0),
	.w3(32'hbbd56512),
	.w4(32'hba067490),
	.w5(32'h3b8b5202),
	.w6(32'hbb858fad),
	.w7(32'h3a8efa43),
	.w8(32'h3b6decd6),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb6dc92),
	.w1(32'hbaf86d14),
	.w2(32'h3b9dae51),
	.w3(32'h3b3d53ef),
	.w4(32'hbb7b7206),
	.w5(32'hb99e424a),
	.w6(32'hbbbd878e),
	.w7(32'hbb71a6eb),
	.w8(32'hba3a4229),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bad6ced),
	.w1(32'h3b0c6e05),
	.w2(32'h3c06ccd8),
	.w3(32'hbb06c0f3),
	.w4(32'hbaf8a8e4),
	.w5(32'h3bc814f8),
	.w6(32'hbbab8a7f),
	.w7(32'hb8d6b0fb),
	.w8(32'h3b25c6da),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b68ebca),
	.w1(32'hbb6035ea),
	.w2(32'hbb0f1820),
	.w3(32'h3b12e6d0),
	.w4(32'hbb252fb7),
	.w5(32'hbb117494),
	.w6(32'hbb056f8b),
	.w7(32'hbb0d0296),
	.w8(32'hbb703d8f),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3958fb69),
	.w1(32'h3b67c38d),
	.w2(32'h3bab60d6),
	.w3(32'hbb54d9c5),
	.w4(32'h3b8ccb4b),
	.w5(32'h3c164a05),
	.w6(32'h3ab960dc),
	.w7(32'h3abb4c57),
	.w8(32'h3c72f066),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c32d723),
	.w1(32'h3bbe65d0),
	.w2(32'h3c057f58),
	.w3(32'h3c64ae8c),
	.w4(32'h3a8ee679),
	.w5(32'h3b67e501),
	.w6(32'hba7c1045),
	.w7(32'h3b38a4d6),
	.w8(32'hbb1fea64),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb39f74d),
	.w1(32'h3b778fe8),
	.w2(32'h3b0e62f8),
	.w3(32'hbbc8c238),
	.w4(32'h3b1e5026),
	.w5(32'h3a2ffb44),
	.w6(32'h3a9fb0de),
	.w7(32'h3aed6fa3),
	.w8(32'h3bb3e220),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb093e9b),
	.w1(32'hbb88d693),
	.w2(32'hbb9306c8),
	.w3(32'hbb3f33f2),
	.w4(32'hbb8527c7),
	.w5(32'hbba429e0),
	.w6(32'hbb47934c),
	.w7(32'hbb83163c),
	.w8(32'hbb83c08f),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9faa83),
	.w1(32'h3b7bd705),
	.w2(32'h3b8ece9c),
	.w3(32'hbba390ce),
	.w4(32'h3adbdc53),
	.w5(32'h3a0b3416),
	.w6(32'h3b442ece),
	.w7(32'h3b687582),
	.w8(32'h3b24c634),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6fd597),
	.w1(32'hbab8205d),
	.w2(32'h3affd5d5),
	.w3(32'hbb109aa0),
	.w4(32'hbb0c5110),
	.w5(32'h3990f588),
	.w6(32'hbb2173dc),
	.w7(32'hbb5abe7f),
	.w8(32'hba45f3e8),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf3b119),
	.w1(32'h3bc32fb0),
	.w2(32'h3c1d4a1f),
	.w3(32'hbb0acfc7),
	.w4(32'h3ab83a1b),
	.w5(32'h3b4c0e42),
	.w6(32'h3b275ccd),
	.w7(32'h3ba157fe),
	.w8(32'h3bd538a3),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b35e980),
	.w1(32'h3822e5fa),
	.w2(32'h39acf59a),
	.w3(32'hbb5fe85d),
	.w4(32'hbb02a2cf),
	.w5(32'hbae5819d),
	.w6(32'hbb89f22b),
	.w7(32'hbb847da2),
	.w8(32'hbb09c6f3),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf7e492),
	.w1(32'hbc06f88d),
	.w2(32'hbc051559),
	.w3(32'hbbe1f178),
	.w4(32'hbbf164e5),
	.w5(32'hbbf39f06),
	.w6(32'hbc036d69),
	.w7(32'hbc08703b),
	.w8(32'hbc003171),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc072daf),
	.w1(32'h3aa086fc),
	.w2(32'h3b5d0ea6),
	.w3(32'hbbfb398d),
	.w4(32'hbb07eb79),
	.w5(32'hba255202),
	.w6(32'hba683eca),
	.w7(32'h3aa08c7c),
	.w8(32'hbab491ab),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa02f8f),
	.w1(32'h3b6a82c9),
	.w2(32'h3ad26fdc),
	.w3(32'hba858e63),
	.w4(32'h3b731cdc),
	.w5(32'h3b0fe77d),
	.w6(32'h3b788225),
	.w7(32'h3b306e9a),
	.w8(32'h3b8c8cbf),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa5a305),
	.w1(32'hbb02b2f3),
	.w2(32'h3b295675),
	.w3(32'h3ab65dae),
	.w4(32'hbb79e5d6),
	.w5(32'hb828639e),
	.w6(32'hbb972571),
	.w7(32'hba7d9e18),
	.w8(32'hbb7f3f0f),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba54cce),
	.w1(32'h3a3dcbbe),
	.w2(32'h3b6310b9),
	.w3(32'hbb67f82c),
	.w4(32'hba91ed54),
	.w5(32'hba698e79),
	.w6(32'hbafa3077),
	.w7(32'h3a9feca5),
	.w8(32'hb96581aa),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7eed474),
	.w1(32'hbc1d88c2),
	.w2(32'hbc018994),
	.w3(32'hbb918833),
	.w4(32'hbc19ae75),
	.w5(32'hbc18943f),
	.w6(32'hbc1d7d76),
	.w7(32'hbc2ecb32),
	.w8(32'hbc2f8b6c),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc08196b),
	.w1(32'h3ba2bc8e),
	.w2(32'h3bd54ca3),
	.w3(32'hbc11662b),
	.w4(32'h3b8f1298),
	.w5(32'h3bb6737e),
	.w6(32'h3bb1905b),
	.w7(32'h3baad7f1),
	.w8(32'h3bde0720),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0e4789),
	.w1(32'h3b9d83b6),
	.w2(32'h3a32834b),
	.w3(32'h3bd784c8),
	.w4(32'h3aebe2f5),
	.w5(32'hba41b297),
	.w6(32'h3b8bbdc7),
	.w7(32'hb88efc48),
	.w8(32'h3ba3bf59),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba494c4a),
	.w1(32'hb9a6f6dd),
	.w2(32'hba9ced47),
	.w3(32'hba8b1f1e),
	.w4(32'h3a07100a),
	.w5(32'hb9e46caa),
	.w6(32'h39872a87),
	.w7(32'hb9fca34a),
	.w8(32'hb992531c),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaf575d),
	.w1(32'h3b299974),
	.w2(32'hb922aa8b),
	.w3(32'hb92246d5),
	.w4(32'hbaf14633),
	.w5(32'hbb2dc90b),
	.w6(32'h3bb0116b),
	.w7(32'h3bc3db10),
	.w8(32'h3bca57e5),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5e49c2),
	.w1(32'h3a91c3db),
	.w2(32'hbadd45fb),
	.w3(32'hba778098),
	.w4(32'h3b3c87f1),
	.w5(32'h39696ba0),
	.w6(32'h3ad2bd52),
	.w7(32'hb9c46b5d),
	.w8(32'h3aec54f8),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396cd09a),
	.w1(32'h3b1aa823),
	.w2(32'h3afd9c24),
	.w3(32'h3b3a7dbb),
	.w4(32'h3b603e5a),
	.w5(32'h3acf9b88),
	.w6(32'h3b0a24eb),
	.w7(32'h3ae78bc8),
	.w8(32'hbb810c11),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9e62ff),
	.w1(32'hba8ff81d),
	.w2(32'hbae3ed6f),
	.w3(32'hbb984c94),
	.w4(32'hba8ce321),
	.w5(32'hbad03a1c),
	.w6(32'h3a90b67c),
	.w7(32'hb9a8b321),
	.w8(32'h393a11d3),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb953d10c),
	.w1(32'h3b26c18c),
	.w2(32'h3b446472),
	.w3(32'hba995308),
	.w4(32'h3b04f363),
	.w5(32'h3af69010),
	.w6(32'hbb01f296),
	.w7(32'hb9821f6e),
	.w8(32'h3abbe0c6),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aace6cd),
	.w1(32'h3b3de72b),
	.w2(32'h3a4661e3),
	.w3(32'hba3d8bb5),
	.w4(32'hba8e5b78),
	.w5(32'hbacf4f4c),
	.w6(32'h39e2b576),
	.w7(32'hbb2b929c),
	.w8(32'h3ba44d19),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2d1ee3),
	.w1(32'hba93a50a),
	.w2(32'hbb0abe77),
	.w3(32'hba84e973),
	.w4(32'hbb8aa749),
	.w5(32'hbbc5955f),
	.w6(32'h3b28c247),
	.w7(32'h37c704c2),
	.w8(32'h3abee209),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdd95eb),
	.w1(32'hbae3d1b4),
	.w2(32'h3be33f68),
	.w3(32'hbc11dffc),
	.w4(32'hbb76bbd1),
	.w5(32'h3ba2f736),
	.w6(32'hbc1235e3),
	.w7(32'hba073eca),
	.w8(32'hbaa03281),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcc2ec0),
	.w1(32'h3b305bec),
	.w2(32'h3b37ef3e),
	.w3(32'h3b6d04bc),
	.w4(32'h394dc57d),
	.w5(32'h3ab5a0ef),
	.w6(32'hbade6d2b),
	.w7(32'h3ab90739),
	.w8(32'h3999e66b),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39faf063),
	.w1(32'h391f759b),
	.w2(32'h3b697f4f),
	.w3(32'hb9ed5a9e),
	.w4(32'hba71a534),
	.w5(32'h3b4985a6),
	.w6(32'hbb575640),
	.w7(32'h3a7d6a06),
	.w8(32'h3a2c80bf),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afeda92),
	.w1(32'hbad6f1fb),
	.w2(32'h3af62637),
	.w3(32'h3a610f15),
	.w4(32'hbaeb607f),
	.w5(32'h3aa674ee),
	.w6(32'hbb85187e),
	.w7(32'hba1436d5),
	.w8(32'hbaa36cbe),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0aae8a),
	.w1(32'hbaa11f52),
	.w2(32'hbae4e3e0),
	.w3(32'hb91fbf29),
	.w4(32'hba17dce1),
	.w5(32'hba9bc12f),
	.w6(32'h38d8c7ff),
	.w7(32'hba0f055d),
	.w8(32'hb9bb1b30),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb084440),
	.w1(32'h3aec9283),
	.w2(32'h3bace7de),
	.w3(32'hbab3db7e),
	.w4(32'hbb480e3f),
	.w5(32'hba5a6db8),
	.w6(32'hbab14f4c),
	.w7(32'h3af978ec),
	.w8(32'hba9f5922),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2ded83),
	.w1(32'hba37397a),
	.w2(32'h3b277ec9),
	.w3(32'hbaaed28a),
	.w4(32'hbaf740e5),
	.w5(32'h3b06a902),
	.w6(32'hbb8084f5),
	.w7(32'hb9769ddb),
	.w8(32'hba1990b1),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3f8469),
	.w1(32'hbc2c5c83),
	.w2(32'hbc273b31),
	.w3(32'h3adf754e),
	.w4(32'hbc2747c9),
	.w5(32'hbc25cf98),
	.w6(32'hbc1b3230),
	.w7(32'hbc21dd09),
	.w8(32'hbc2109fc),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3708b0),
	.w1(32'hbad397da),
	.w2(32'h3bb08358),
	.w3(32'hbc27dd06),
	.w4(32'hbae405a7),
	.w5(32'h3b9de294),
	.w6(32'hbb2f989f),
	.w7(32'h3ab692e3),
	.w8(32'h3ad8c369),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf8a22d),
	.w1(32'hbb0229e4),
	.w2(32'h3bf45e51),
	.w3(32'h3b8780d3),
	.w4(32'hbb4ccd1d),
	.w5(32'h3bd746e8),
	.w6(32'hbbb77c2b),
	.w7(32'h3bdf5375),
	.w8(32'h3a6651dc),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a7691),
	.w1(32'h3b85ba65),
	.w2(32'h3c0bc699),
	.w3(32'hbb99e6e4),
	.w4(32'h3b0fcf5f),
	.w5(32'h3bd73d3f),
	.w6(32'hbada0e96),
	.w7(32'h3b874a8a),
	.w8(32'h3b813832),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcb1013),
	.w1(32'hbb1bec75),
	.w2(32'hbb34688c),
	.w3(32'h3b89a509),
	.w4(32'hbb31df28),
	.w5(32'hbb4ee78b),
	.w6(32'hbb5917e9),
	.w7(32'hbb451111),
	.w8(32'hbb0cdf41),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a4bf4),
	.w1(32'hbaa74f9d),
	.w2(32'h3b863ec9),
	.w3(32'hbb86cc8f),
	.w4(32'hbb362709),
	.w5(32'h3b40c209),
	.w6(32'hba189782),
	.w7(32'h3ae42ebf),
	.w8(32'h3a946be0),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7c8727),
	.w1(32'hba60a34f),
	.w2(32'h3b86e086),
	.w3(32'h3ae1edf4),
	.w4(32'hbb2528fb),
	.w5(32'h3b5e7e76),
	.w6(32'hbbaf83e9),
	.w7(32'h38b6d2d6),
	.w8(32'hb9a97f54),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9da6dc),
	.w1(32'h3a84d6de),
	.w2(32'h3b40f67a),
	.w3(32'h3b4424aa),
	.w4(32'hba918c59),
	.w5(32'h3ac736fd),
	.w6(32'hba6ec90c),
	.w7(32'h3b0abe78),
	.w8(32'h3a65a03e),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3fd2d6),
	.w1(32'h3b11d424),
	.w2(32'h3b9c4f28),
	.w3(32'h3a9e23a8),
	.w4(32'hb6e4367e),
	.w5(32'h3b5f0c88),
	.w6(32'hba02402d),
	.w7(32'h3b4b8c5f),
	.w8(32'h3af47af9),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba99beb),
	.w1(32'hbaf57146),
	.w2(32'h39f71ba3),
	.w3(32'h3b280319),
	.w4(32'hbbbd187a),
	.w5(32'hbb9211dd),
	.w6(32'hba89867b),
	.w7(32'h3b3210c6),
	.w8(32'hb9274bf1),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38db3ac0),
	.w1(32'h3a552bd3),
	.w2(32'hbb4c6472),
	.w3(32'hbbb3a4db),
	.w4(32'h39fca296),
	.w5(32'hbb4ef1e4),
	.w6(32'h3aa245e8),
	.w7(32'hbb26b214),
	.w8(32'h3ad4bf8c),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ae7d1f),
	.w1(32'h3b388549),
	.w2(32'h39bea23d),
	.w3(32'h3a4c26bf),
	.w4(32'h3a31bd30),
	.w5(32'hba37f6e2),
	.w6(32'h3a985a0b),
	.w7(32'hb9f4b252),
	.w8(32'hbb08d359),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398ad412),
	.w1(32'h38f0bb44),
	.w2(32'h3abc9b20),
	.w3(32'hbaa6a8d9),
	.w4(32'hba8f074e),
	.w5(32'h39c8843c),
	.w6(32'h3989c981),
	.w7(32'h3b1a034f),
	.w8(32'hbb02115b),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8ca54b),
	.w1(32'hb9d08b4d),
	.w2(32'h3b24b09d),
	.w3(32'hbab0e95c),
	.w4(32'hbaeb02e2),
	.w5(32'h3aeefe97),
	.w6(32'hbb3b322f),
	.w7(32'h3a6fac0c),
	.w8(32'hba43edf5),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b04482d),
	.w1(32'hbb7f5b7c),
	.w2(32'hbb2e5d08),
	.w3(32'h394f96ac),
	.w4(32'hbbe8a585),
	.w5(32'hbbd71762),
	.w6(32'hbaadf74a),
	.w7(32'h3a43e92f),
	.w8(32'hb8cdf2a1),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf12c64),
	.w1(32'h3c15366b),
	.w2(32'h3c0d99f7),
	.w3(32'hbbdc737e),
	.w4(32'h3bcc6081),
	.w5(32'h3bda78c1),
	.w6(32'h3c0c5d58),
	.w7(32'h3c28a505),
	.w8(32'h3c2919cf),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3b588b),
	.w1(32'h3c1172e7),
	.w2(32'h3c1662ca),
	.w3(32'h3c1283f5),
	.w4(32'h3ab86bc5),
	.w5(32'h3af74b81),
	.w6(32'h3b5bdbfe),
	.w7(32'h3b9e0113),
	.w8(32'hbb0e5674),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6719b9),
	.w1(32'hb9a3da9a),
	.w2(32'hb9da3446),
	.w3(32'hbb100114),
	.w4(32'hb9b44614),
	.w5(32'hb9bcdbd5),
	.w6(32'hb992df82),
	.w7(32'hb994632f),
	.w8(32'hb9520f16),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab80039),
	.w1(32'h3a9d676f),
	.w2(32'h3ac49ec6),
	.w3(32'h3af10c08),
	.w4(32'h3994d80d),
	.w5(32'hba27ed89),
	.w6(32'h3b216bd0),
	.w7(32'h3a5660b2),
	.w8(32'h39dbd7b1),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule