module layer_8_featuremap_57(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b532ce),
	.w1(32'hb9f3c22e),
	.w2(32'hba7b6cf4),
	.w3(32'h3a1f34c2),
	.w4(32'hba250dde),
	.w5(32'hb950c5a0),
	.w6(32'hba424b3f),
	.w7(32'hba57f4e9),
	.w8(32'hba71cad3),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38090dbf),
	.w1(32'h392c192c),
	.w2(32'hb9703aaa),
	.w3(32'h38e2f24c),
	.w4(32'hb895a3ac),
	.w5(32'h37f5e4e7),
	.w6(32'hb90b7c37),
	.w7(32'hb8ca6519),
	.w8(32'hba3469d1),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb78c5c60),
	.w1(32'h393c301a),
	.w2(32'hb8d7757b),
	.w3(32'h383e6eac),
	.w4(32'hb92b9d9d),
	.w5(32'hb915f4de),
	.w6(32'hb913a1a2),
	.w7(32'hb8c519dc),
	.w8(32'hba288780),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacf248b),
	.w1(32'hbaed4810),
	.w2(32'hbacb28e4),
	.w3(32'hba9ee6a5),
	.w4(32'hba16e2ad),
	.w5(32'hbaa0f72b),
	.w6(32'hb9a0b5c7),
	.w7(32'hba720f60),
	.w8(32'hba67ff83),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ec8be4),
	.w1(32'h39eddff5),
	.w2(32'h38fc810a),
	.w3(32'h3a1d5410),
	.w4(32'h3996294f),
	.w5(32'hb9602f7f),
	.w6(32'h39a505d4),
	.w7(32'h39bf2552),
	.w8(32'hbaa682ac),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba36ed82),
	.w1(32'h391c731a),
	.w2(32'h3a6007c8),
	.w3(32'hb896f036),
	.w4(32'h39102360),
	.w5(32'h3a81ffb2),
	.w6(32'hb9feb8e1),
	.w7(32'h3aad465b),
	.w8(32'hb98cde1e),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h370f6863),
	.w1(32'h38867cf8),
	.w2(32'hba069de6),
	.w3(32'h39221ca6),
	.w4(32'hb9f8762b),
	.w5(32'hba2617b1),
	.w6(32'hb956c575),
	.w7(32'hb8c43e2c),
	.w8(32'hb9e5f7ca),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8ea89a),
	.w1(32'h3a89fba3),
	.w2(32'h3a06f80b),
	.w3(32'h3a5e0d04),
	.w4(32'h3a01ae9a),
	.w5(32'hb88cd840),
	.w6(32'h3a731d76),
	.w7(32'h3a74795e),
	.w8(32'hba41e027),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h396f4b37),
	.w1(32'h38abd0c2),
	.w2(32'hb9c1dcdf),
	.w3(32'h3a1dd557),
	.w4(32'hb94b3541),
	.w5(32'hb9ce730d),
	.w6(32'hb97cddbb),
	.w7(32'hb9930e0c),
	.w8(32'hb8f8d321),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab75cc6),
	.w1(32'hbae6a579),
	.w2(32'hb96708f1),
	.w3(32'h39276ac0),
	.w4(32'h3a9ca148),
	.w5(32'hb69346e1),
	.w6(32'h3a233dba),
	.w7(32'hbad85183),
	.w8(32'hbaceb347),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3d05b5),
	.w1(32'hb9f1d70d),
	.w2(32'hbaa979b5),
	.w3(32'hba79ab7c),
	.w4(32'hba8fd666),
	.w5(32'hbaa7b20b),
	.w6(32'hba9e57ac),
	.w7(32'hba335be6),
	.w8(32'hba9417a0),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4454a2),
	.w1(32'hb987cced),
	.w2(32'hba8a43ab),
	.w3(32'hb955ad89),
	.w4(32'hb959aa76),
	.w5(32'hb9b43394),
	.w6(32'hba80fe60),
	.w7(32'hb98ab3f3),
	.w8(32'hba39116c),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e75147),
	.w1(32'h38af3034),
	.w2(32'hba0bef8b),
	.w3(32'hb8ef7dcf),
	.w4(32'hb8101bcf),
	.w5(32'hb9a4aef1),
	.w6(32'hb982a9a4),
	.w7(32'h38edbbd9),
	.w8(32'hbaaa515c),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92d146e),
	.w1(32'hba079692),
	.w2(32'h39d8a38a),
	.w3(32'h39ba8855),
	.w4(32'hba91aaaa),
	.w5(32'h3a594e41),
	.w6(32'hba1bcd59),
	.w7(32'h39a76171),
	.w8(32'hba8b3bb5),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8cf48b0),
	.w1(32'hb9690752),
	.w2(32'h396aa332),
	.w3(32'h39a15912),
	.w4(32'hb9e4eac1),
	.w5(32'h3922a0f1),
	.w6(32'hb911c163),
	.w7(32'h38df7199),
	.w8(32'h39972cc7),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c2c3ad),
	.w1(32'h387fb3bd),
	.w2(32'hb8a5618a),
	.w3(32'h396cb991),
	.w4(32'hba6c794c),
	.w5(32'hb98928df),
	.w6(32'h39174156),
	.w7(32'hb90ee2f5),
	.w8(32'hb9156fe6),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac3e514),
	.w1(32'hb99c9686),
	.w2(32'hb96413ab),
	.w3(32'hbac43656),
	.w4(32'h3a0233ab),
	.w5(32'h3a00d808),
	.w6(32'hbaca038e),
	.w7(32'hbb3fb4e5),
	.w8(32'hbacaa2f6),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba88f25e),
	.w1(32'hb7b3611a),
	.w2(32'hb9bb293c),
	.w3(32'hb9f80371),
	.w4(32'hba054194),
	.w5(32'hb9bafe48),
	.w6(32'hba5aa463),
	.w7(32'hb9d10210),
	.w8(32'hb990b78b),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e96feb),
	.w1(32'hbaf8853a),
	.w2(32'hbb5b081c),
	.w3(32'hbaf476ce),
	.w4(32'hbb3d5894),
	.w5(32'hbb544f9a),
	.w6(32'hbb437144),
	.w7(32'hbb157e56),
	.w8(32'hbba4e328),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7f82f2),
	.w1(32'h3bd99d9b),
	.w2(32'hbb0c3367),
	.w3(32'hbb0cd0a5),
	.w4(32'h3a971d6c),
	.w5(32'hbb07db70),
	.w6(32'h39ac02f6),
	.w7(32'h3aa731c7),
	.w8(32'hba3ea22d),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba951ead),
	.w1(32'hb93753fd),
	.w2(32'h397e4ee5),
	.w3(32'h3927d46d),
	.w4(32'h3a07a59d),
	.w5(32'hb96545f1),
	.w6(32'hba841bec),
	.w7(32'hb9b62958),
	.w8(32'hba388714),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1fdf8b),
	.w1(32'h3a534562),
	.w2(32'h39bfd27f),
	.w3(32'h3a101f16),
	.w4(32'h38adaa42),
	.w5(32'hb989c2bc),
	.w6(32'h38aba899),
	.w7(32'h3a10cea7),
	.w8(32'h3b3c7aae),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad4c4bd),
	.w1(32'hb9c2122c),
	.w2(32'hba4874a6),
	.w3(32'h39ab8deb),
	.w4(32'h3976cc6b),
	.w5(32'h3a69c506),
	.w6(32'hb9449148),
	.w7(32'h3a198b40),
	.w8(32'hbab3169e),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb87bebe4),
	.w1(32'hb903a03d),
	.w2(32'hb8dd65c2),
	.w3(32'h38995642),
	.w4(32'hb9e67628),
	.w5(32'h39b49795),
	.w6(32'hba594325),
	.w7(32'hb976a6bd),
	.w8(32'h38232fb3),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba53fe6c),
	.w1(32'h397eae42),
	.w2(32'hba45e7a2),
	.w3(32'hbb0936f7),
	.w4(32'hba920f51),
	.w5(32'hba9783ac),
	.w6(32'hba707622),
	.w7(32'hba8b5756),
	.w8(32'h3b3322bb),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a309db6),
	.w1(32'hb911f948),
	.w2(32'h3988bf89),
	.w3(32'h3a3688b7),
	.w4(32'h39fd38c1),
	.w5(32'h3a155f8a),
	.w6(32'h39a6c563),
	.w7(32'h3ac7eacf),
	.w8(32'h3b15089d),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab1b64a),
	.w1(32'h398305aa),
	.w2(32'h3a794a24),
	.w3(32'h3a8b2c0c),
	.w4(32'h3a41088a),
	.w5(32'h3a61d04d),
	.w6(32'h39c5f95e),
	.w7(32'h3a99688d),
	.w8(32'hb9b8e64b),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1c4227),
	.w1(32'h3bec3ab4),
	.w2(32'h3bb01716),
	.w3(32'hbb86a210),
	.w4(32'h3a238d54),
	.w5(32'hbb4a001f),
	.w6(32'hbb2c0dd6),
	.w7(32'h39fd3658),
	.w8(32'h3c1a8867),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1347ac),
	.w1(32'hbaa440d0),
	.w2(32'hbaa6df3b),
	.w3(32'hb90d7c81),
	.w4(32'hbb45c75a),
	.w5(32'hba80ccb7),
	.w6(32'h3985108c),
	.w7(32'hbb054fa3),
	.w8(32'hba997370),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b3a4d9),
	.w1(32'hb91a3ebb),
	.w2(32'hb995c98c),
	.w3(32'hb9056cf8),
	.w4(32'hb915f2b6),
	.w5(32'hb96067da),
	.w6(32'hb9bb748a),
	.w7(32'hb9465fa5),
	.w8(32'hbb0b1ed1),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1d3f6f),
	.w1(32'h3b06792b),
	.w2(32'hba73570c),
	.w3(32'hbb19f2ab),
	.w4(32'h3abe27c6),
	.w5(32'hb91d2d48),
	.w6(32'hbb17b8f9),
	.w7(32'hba4c9746),
	.w8(32'hba2b71cf),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8d12c2),
	.w1(32'hba550a1f),
	.w2(32'h3983816e),
	.w3(32'hb936fa3f),
	.w4(32'hba1393c5),
	.w5(32'hba858f25),
	.w6(32'hbaa72397),
	.w7(32'h3a65fc77),
	.w8(32'hbafafd1c),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb39d0ab),
	.w1(32'hbaf44370),
	.w2(32'hba851b48),
	.w3(32'hbb010077),
	.w4(32'h39dc1e3d),
	.w5(32'h3a2c493c),
	.w6(32'hb99cc603),
	.w7(32'hb9dbf1b8),
	.w8(32'hbb157265),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab583d7),
	.w1(32'h3b8ddc5b),
	.w2(32'h3a91f327),
	.w3(32'hbab2214c),
	.w4(32'hba44cd3b),
	.w5(32'h3b03431f),
	.w6(32'hbb1c6057),
	.w7(32'hba147787),
	.w8(32'hba8756fd),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac253b4),
	.w1(32'hba17e6d9),
	.w2(32'h395ff948),
	.w3(32'hba483bfa),
	.w4(32'hba632b6f),
	.w5(32'h3a1876d1),
	.w6(32'hbae63d5f),
	.w7(32'h3893caf2),
	.w8(32'hba3fa4ef),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4b9d3c),
	.w1(32'h39991077),
	.w2(32'hb9d72de3),
	.w3(32'h38edf53d),
	.w4(32'hbabf9254),
	.w5(32'hb8d16673),
	.w6(32'hba16015b),
	.w7(32'hb9fede0c),
	.w8(32'hbaad59c9),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394933eb),
	.w1(32'hb9a1acba),
	.w2(32'hba3954b1),
	.w3(32'hba8b45d9),
	.w4(32'hba5f92a2),
	.w5(32'h3721ab5c),
	.w6(32'hbaae7d19),
	.w7(32'hba6541c9),
	.w8(32'hba6b9e16),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8516e74),
	.w1(32'hb8b13746),
	.w2(32'hb9da287e),
	.w3(32'h39020175),
	.w4(32'hb99e3790),
	.w5(32'hba006de9),
	.w6(32'hb943b379),
	.w7(32'hb965de91),
	.w8(32'hbaf659f4),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h381dfdf1),
	.w1(32'hb94269f0),
	.w2(32'h3a3e2ccb),
	.w3(32'h3a58ca64),
	.w4(32'hba0c69e0),
	.w5(32'h398e1359),
	.w6(32'h37cff985),
	.w7(32'h39ece7e6),
	.w8(32'hba4bc4d7),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99d357c),
	.w1(32'hb9c6bca3),
	.w2(32'hba02eb1d),
	.w3(32'hba496d78),
	.w4(32'hba9f23bb),
	.w5(32'hba812163),
	.w6(32'hba342ccc),
	.w7(32'hb954f0f3),
	.w8(32'h3a92a1c7),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0834f8),
	.w1(32'hba20f74f),
	.w2(32'hba0d4574),
	.w3(32'hbadf330e),
	.w4(32'h39adcebc),
	.w5(32'h3a88aef9),
	.w6(32'hbb42ce28),
	.w7(32'h3a0b2fdc),
	.w8(32'h3b4a9ea8),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb32eeee),
	.w1(32'hbb309de5),
	.w2(32'hba59ea87),
	.w3(32'h3bca1a93),
	.w4(32'h3b0929f0),
	.w5(32'hbad74d68),
	.w6(32'h3a029efd),
	.w7(32'hba25f3bd),
	.w8(32'hbb6914cf),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafb5ac8),
	.w1(32'h3c9cc705),
	.w2(32'hbbe02140),
	.w3(32'h3b9fa7a1),
	.w4(32'h3b884889),
	.w5(32'hbbe4c6a5),
	.w6(32'hba422749),
	.w7(32'hbbd6f3ae),
	.w8(32'h3a0171e3),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc151e0d),
	.w1(32'hbbd3c2a7),
	.w2(32'h3bb1e1f7),
	.w3(32'hbb5cab56),
	.w4(32'hbbc84e50),
	.w5(32'hb83ac99d),
	.w6(32'hbb9e0d85),
	.w7(32'h3b3bc16a),
	.w8(32'h3ac90817),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad88371),
	.w1(32'hbc13201f),
	.w2(32'hbc83b0d6),
	.w3(32'h3ad74a04),
	.w4(32'hbbf8897d),
	.w5(32'hbc801426),
	.w6(32'hbc10b417),
	.w7(32'hbc832123),
	.w8(32'h3c408ad4),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c404e0c),
	.w1(32'h3a308211),
	.w2(32'hbc73510d),
	.w3(32'h3c70f488),
	.w4(32'h3baf43ab),
	.w5(32'hbb9e5e89),
	.w6(32'h3b75eb12),
	.w7(32'hbc6242ee),
	.w8(32'h3bc26528),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaed434),
	.w1(32'h3baeb733),
	.w2(32'hb99f7903),
	.w3(32'hbc420ae2),
	.w4(32'h3ba7c535),
	.w5(32'h3bd87518),
	.w6(32'h3bc683cf),
	.w7(32'hbcf53dd8),
	.w8(32'h3bd1784c),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2e324e),
	.w1(32'hbc04dbda),
	.w2(32'hbcb22181),
	.w3(32'h3c8b38bc),
	.w4(32'hb918c4d0),
	.w5(32'hbc5f1a87),
	.w6(32'hbc5fca0f),
	.w7(32'hbc241413),
	.w8(32'h3c4a781e),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d1c9699),
	.w1(32'h3b9abc17),
	.w2(32'hbc800bf0),
	.w3(32'h3ca9a61a),
	.w4(32'h3b8119d1),
	.w5(32'hbbc4c479),
	.w6(32'hbbae706f),
	.w7(32'hbc097ca5),
	.w8(32'h3ba4b44e),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a679c38),
	.w1(32'hbbf2ddf1),
	.w2(32'hbc3b9093),
	.w3(32'h3bba65f3),
	.w4(32'hbb8c6053),
	.w5(32'hbc387972),
	.w6(32'hbbf4b451),
	.w7(32'hbc62cc5e),
	.w8(32'hbaf43d98),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeb1613),
	.w1(32'h3a19db5f),
	.w2(32'h3b2d4c40),
	.w3(32'hbb3ea8cf),
	.w4(32'h3a41ac2d),
	.w5(32'h3a4f59fe),
	.w6(32'h3adfe20e),
	.w7(32'h3b09e007),
	.w8(32'hbb239132),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc85f2ed),
	.w1(32'hbaeffd22),
	.w2(32'h3b8b1b4a),
	.w3(32'hbc113fbf),
	.w4(32'hbb08c951),
	.w5(32'hbb123c32),
	.w6(32'h3b11a22f),
	.w7(32'h3b8726b2),
	.w8(32'hbc34ca23),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd0d1d8),
	.w1(32'hbc969bd3),
	.w2(32'h3c2de8a9),
	.w3(32'hbca033e2),
	.w4(32'hbcc4be01),
	.w5(32'hbb1851c6),
	.w6(32'hbc917c16),
	.w7(32'hbc104f65),
	.w8(32'h3d1dbea2),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d69cd10),
	.w1(32'h3c54f640),
	.w2(32'hbd251a82),
	.w3(32'h3d44d0a1),
	.w4(32'h3ca62bd9),
	.w5(32'hbca57437),
	.w6(32'h3ad66522),
	.w7(32'hbd1f332b),
	.w8(32'hbc487e85),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a2420a),
	.w1(32'h3c2210c8),
	.w2(32'hba7de4b8),
	.w3(32'hbba139b0),
	.w4(32'hbaa8fc79),
	.w5(32'h3b41ccf5),
	.w6(32'hbc381f2b),
	.w7(32'hbc89206d),
	.w8(32'h3c676205),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf22091),
	.w1(32'hba47cf36),
	.w2(32'h3c552879),
	.w3(32'h3c00a267),
	.w4(32'h3b9e17b0),
	.w5(32'hbb266c57),
	.w6(32'h3bbd43c9),
	.w7(32'h3be442fb),
	.w8(32'h3c148bdd),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8ad272),
	.w1(32'hbca4fafc),
	.w2(32'hbbd40006),
	.w3(32'hbb5f066a),
	.w4(32'hbc96ea8c),
	.w5(32'h3ba147ba),
	.w6(32'hbcb80479),
	.w7(32'hbb6d62cd),
	.w8(32'hbc16f765),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba629ba3),
	.w1(32'hbb8c1288),
	.w2(32'h3b986989),
	.w3(32'hbba02e48),
	.w4(32'h3bac7552),
	.w5(32'hbc04b082),
	.w6(32'hbb507a92),
	.w7(32'hba0a44dc),
	.w8(32'hbc58593d),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc619cd1),
	.w1(32'hba7b6d14),
	.w2(32'h3ccb1fbb),
	.w3(32'hbc9581b1),
	.w4(32'hbc22f5d7),
	.w5(32'h3c3d8e5f),
	.w6(32'hbbab8764),
	.w7(32'h3ca6c532),
	.w8(32'h3ace063e),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c47323a),
	.w1(32'hbb767971),
	.w2(32'hbc81bf64),
	.w3(32'h3b4bd115),
	.w4(32'hbb9c9e36),
	.w5(32'h3b2e148b),
	.w6(32'hbc53995b),
	.w7(32'hbc10ff1c),
	.w8(32'hbc036244),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2f6acf),
	.w1(32'h3cb69bbf),
	.w2(32'hbbc73973),
	.w3(32'hbcf71c8b),
	.w4(32'hbc2b1741),
	.w5(32'h3bd54d16),
	.w6(32'hbb0e0802),
	.w7(32'hbbd55ca0),
	.w8(32'h3c6c4324),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbdc646),
	.w1(32'hbaa1d3ea),
	.w2(32'hbc0811cd),
	.w3(32'h3c744afe),
	.w4(32'h3c017ece),
	.w5(32'hbb0d25f1),
	.w6(32'hba069e48),
	.w7(32'hbbd48867),
	.w8(32'h3ae8adbb),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb97b525),
	.w1(32'h397caace),
	.w2(32'hbc1b78c8),
	.w3(32'hb915e8a4),
	.w4(32'h3b002433),
	.w5(32'hbc1457aa),
	.w6(32'hbaab448e),
	.w7(32'hbc4c1c04),
	.w8(32'hbccae6a0),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc12851f),
	.w1(32'h3c4de5e2),
	.w2(32'hbb89c58f),
	.w3(32'hbabe8a50),
	.w4(32'h3a0dfa17),
	.w5(32'hbc259931),
	.w6(32'hbb009cb2),
	.w7(32'h3c2672de),
	.w8(32'h3b86cc1f),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92a69bb),
	.w1(32'hbc0f5d8d),
	.w2(32'hbb031dd9),
	.w3(32'h3b308104),
	.w4(32'hbc316403),
	.w5(32'hbb611773),
	.w6(32'hbc191ba1),
	.w7(32'hbb42046f),
	.w8(32'hb858e840),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f97d4),
	.w1(32'hba035a5d),
	.w2(32'h3ba36b34),
	.w3(32'hbae77fa5),
	.w4(32'hba938509),
	.w5(32'h3aa75c65),
	.w6(32'h398c350f),
	.w7(32'h3b263ff9),
	.w8(32'hba4edff5),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba74f31),
	.w1(32'h397602c7),
	.w2(32'h39fa2c83),
	.w3(32'hbb145091),
	.w4(32'hb8560f3e),
	.w5(32'hba4241b7),
	.w6(32'h3a8845ec),
	.w7(32'h39b45455),
	.w8(32'h3c27373f),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc7d6520),
	.w1(32'hbbffc30c),
	.w2(32'hbc0ca105),
	.w3(32'hbae18fb1),
	.w4(32'h3b36c4f4),
	.w5(32'h3b2591b5),
	.w6(32'hbbc28468),
	.w7(32'hbc009196),
	.w8(32'h3b7809be),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c99ff1),
	.w1(32'hbba46b7a),
	.w2(32'hbc3684c0),
	.w3(32'h3bb9668d),
	.w4(32'hbb114c9d),
	.w5(32'hbc0f6524),
	.w6(32'hbbabee41),
	.w7(32'hbc55a0d1),
	.w8(32'hbd144719),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd84647b),
	.w1(32'hbbbded99),
	.w2(32'h3d6f26d6),
	.w3(32'hbd5c0196),
	.w4(32'hbcaea582),
	.w5(32'h3cd9019d),
	.w6(32'hbb3c61f1),
	.w7(32'h3d28ee98),
	.w8(32'h3aa27c27),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3d5078),
	.w1(32'hbb100e25),
	.w2(32'hb99467ea),
	.w3(32'h3b1fb2a3),
	.w4(32'hba2005e7),
	.w5(32'hbb1c31c5),
	.w6(32'hb801c1cc),
	.w7(32'hba513270),
	.w8(32'h3bb7a439),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5af6c7),
	.w1(32'hbbaaa709),
	.w2(32'hbc30e10a),
	.w3(32'h3c1681d0),
	.w4(32'hb96e097e),
	.w5(32'hbc010161),
	.w6(32'hbbbbf2fb),
	.w7(32'hbc509f70),
	.w8(32'h3ac483a2),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb88953e),
	.w1(32'hbae2cca8),
	.w2(32'hba2f9772),
	.w3(32'h3acd47b9),
	.w4(32'hb8d4784e),
	.w5(32'hbb400c83),
	.w6(32'h3a040aff),
	.w7(32'hbb1a849e),
	.w8(32'h3bfb5b71),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9f8596),
	.w1(32'hbcccc694),
	.w2(32'hbc6c4efc),
	.w3(32'h3b73f23f),
	.w4(32'h3b8b09ee),
	.w5(32'h3bd998d1),
	.w6(32'h3c75e9f4),
	.w7(32'h3b7b42ff),
	.w8(32'h3b81327d),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad36030),
	.w1(32'hba7bfe0d),
	.w2(32'hbc0ebf9b),
	.w3(32'h3c0197d9),
	.w4(32'h3b69150f),
	.w5(32'hbb7bb383),
	.w6(32'h3ab62029),
	.w7(32'hbbe528b8),
	.w8(32'h374fa990),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb35851),
	.w1(32'hba89d3bd),
	.w2(32'h3b445344),
	.w3(32'hb9b6ec71),
	.w4(32'hb992a776),
	.w5(32'hb9fdb1f7),
	.w6(32'h399fcd06),
	.w7(32'h3aa07a15),
	.w8(32'h3aa6c0f8),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7d0400),
	.w1(32'hbb2a03cd),
	.w2(32'hbb954284),
	.w3(32'h3b87d805),
	.w4(32'h3b0060f0),
	.w5(32'hbb319138),
	.w6(32'hb9b04c9d),
	.w7(32'hbb3e6faf),
	.w8(32'hbd2c9141),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd951c2d),
	.w1(32'hbbdc3a05),
	.w2(32'h3d8e8d16),
	.w3(32'hbd7be66f),
	.w4(32'hbcc07243),
	.w5(32'h3d0592eb),
	.w6(32'hbb6d8480),
	.w7(32'h3d4e3baf),
	.w8(32'hbc853d49),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd0f99cc),
	.w1(32'hbb49040d),
	.w2(32'h3d02e705),
	.w3(32'hbcccc5c1),
	.w4(32'hbbdaa889),
	.w5(32'h3c7631e2),
	.w6(32'h3b2745f2),
	.w7(32'h3cad47ab),
	.w8(32'h3b24b49b),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb206d60),
	.w1(32'hbc2bedb6),
	.w2(32'h3b4961f0),
	.w3(32'h3ad3128c),
	.w4(32'hbc2615e4),
	.w5(32'h3a082f39),
	.w6(32'hbc31829e),
	.w7(32'h3a461615),
	.w8(32'h3b766573),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b208cc1),
	.w1(32'h39c67024),
	.w2(32'hbc8d0525),
	.w3(32'hbcbae0bb),
	.w4(32'hbc2e8d40),
	.w5(32'h3bb93ab8),
	.w6(32'hba3455dd),
	.w7(32'hba40bd20),
	.w8(32'h3bbddaed),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb926f4ac),
	.w1(32'h3a2da0c8),
	.w2(32'hbbe8bc81),
	.w3(32'h3bbb10c6),
	.w4(32'h3b015091),
	.w5(32'hbb5d1a56),
	.w6(32'h3b35fc17),
	.w7(32'hbba5c87e),
	.w8(32'h3c3d226c),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bacda95),
	.w1(32'hbc52ec22),
	.w2(32'hbc947d53),
	.w3(32'h3c746562),
	.w4(32'hbb40bb9a),
	.w5(32'hbc577a8a),
	.w6(32'hbc3d3617),
	.w7(32'hbc9d7052),
	.w8(32'hbb332c7f),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbde9a9),
	.w1(32'hbc8aebab),
	.w2(32'hbb769bf9),
	.w3(32'hbc3e34de),
	.w4(32'hbc2542c6),
	.w5(32'h3bba33c0),
	.w6(32'hbd062566),
	.w7(32'hbbf6b6ff),
	.w8(32'h3cadd005),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d199c1d),
	.w1(32'h3ba162c7),
	.w2(32'hbd04eff7),
	.w3(32'h3d09f174),
	.w4(32'h3c36abe4),
	.w5(32'hbc92eee5),
	.w6(32'hbbfbd211),
	.w7(32'hbd04d6c5),
	.w8(32'h3b2daf08),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2dc3f3),
	.w1(32'hbbc40d48),
	.w2(32'hbc4df7b3),
	.w3(32'h3b867e69),
	.w4(32'hbb2d5d2d),
	.w5(32'hbc391c0d),
	.w6(32'hbbcfd744),
	.w7(32'hbc65ee24),
	.w8(32'h3c7e7edc),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d520857),
	.w1(32'h3bca7981),
	.w2(32'hbca76c1e),
	.w3(32'h3ce3f962),
	.w4(32'h3ba72571),
	.w5(32'hbc016f92),
	.w6(32'hbbd84b22),
	.w7(32'hbc351b6b),
	.w8(32'h3c170fd4),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be2d37e),
	.w1(32'hbc080a68),
	.w2(32'hbc891610),
	.w3(32'h3c1e0f5c),
	.w4(32'hbc2faa7c),
	.w5(32'hbc76eb51),
	.w6(32'hbc20af15),
	.w7(32'hbc75e90d),
	.w8(32'h3bf84742),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cdbb3e2),
	.w1(32'h3b9a7b54),
	.w2(32'hbce25799),
	.w3(32'h3ca2169a),
	.w4(32'h3c0e8f22),
	.w5(32'hbc35a5e7),
	.w6(32'hbba71cc0),
	.w7(32'hbc6ccf24),
	.w8(32'h3c832490),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d447023),
	.w1(32'h3bbd7fa4),
	.w2(32'hbc9cb39d),
	.w3(32'h3cd61914),
	.w4(32'h3b9e725a),
	.w5(32'hbbef0517),
	.w6(32'hbbc96884),
	.w7(32'hbc29e017),
	.w8(32'h3c61b081),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d247382),
	.w1(32'h3b9556d4),
	.w2(32'hbc89ed6e),
	.w3(32'h3cb33476),
	.w4(32'h3b860fe4),
	.w5(32'hbbd91178),
	.w6(32'hbbbcf9f2),
	.w7(32'hbc154002),
	.w8(32'h3cdc5336),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d334ce3),
	.w1(32'h3bd481a7),
	.w2(32'hbd160cd4),
	.w3(32'h3d15b119),
	.w4(32'h3c5a0f3c),
	.w5(32'hbca54b77),
	.w6(32'hbb2072ed),
	.w7(32'hbd11e5ac),
	.w8(32'hba53e1ad),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b03b38e),
	.w1(32'hbd2ba852),
	.w2(32'hbc1b6979),
	.w3(32'hbabd957d),
	.w4(32'hbd64db02),
	.w5(32'hbc49d7ff),
	.w6(32'hbd5b62a5),
	.w7(32'hbcafff26),
	.w8(32'hbab61490),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc2c61f),
	.w1(32'hba541a01),
	.w2(32'h3ad50d89),
	.w3(32'hbb3de4cf),
	.w4(32'hb9829f6b),
	.w5(32'h398f2c1c),
	.w6(32'h3a3768ea),
	.w7(32'h3ab86549),
	.w8(32'hbb8a45bd),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a45805c),
	.w1(32'hbbe71db8),
	.w2(32'hbba4df01),
	.w3(32'h3ceab6f7),
	.w4(32'h3c06f709),
	.w5(32'hbc6a751e),
	.w6(32'h3b7fdeeb),
	.w7(32'h3c4929d2),
	.w8(32'h3cf93194),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d6bb9b7),
	.w1(32'h3b840142),
	.w2(32'hbd6febda),
	.w3(32'h3d4ff299),
	.w4(32'h3c73b519),
	.w5(32'hbd060526),
	.w6(32'hbc1d75e7),
	.w7(32'hbd4396fc),
	.w8(32'h3b2839b3),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8089c1),
	.w1(32'hbbcb443a),
	.w2(32'hba8b0b09),
	.w3(32'h3c8bae2c),
	.w4(32'h3af21e28),
	.w5(32'hbc41127d),
	.w6(32'hbc1c79cc),
	.w7(32'hbc528410),
	.w8(32'h3a7b7565),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5e2b69),
	.w1(32'h3c50281f),
	.w2(32'hbb56b74e),
	.w3(32'hba94f607),
	.w4(32'h3aef4ff3),
	.w5(32'h39ceea90),
	.w6(32'h3be0c6c3),
	.w7(32'hbaab667c),
	.w8(32'hbd172dd1),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd8161ab),
	.w1(32'hbbb5aa21),
	.w2(32'h3d7e16a5),
	.w3(32'hbd58baf0),
	.w4(32'hbca3e619),
	.w5(32'h3cf17975),
	.w6(32'hbb0a91d0),
	.w7(32'h3d360533),
	.w8(32'h3c1639bb),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1e1062),
	.w1(32'hbbe7061e),
	.w2(32'hbbbb588d),
	.w3(32'h3bcf4e8f),
	.w4(32'hbbe5a566),
	.w5(32'hbbff7348),
	.w6(32'hbc053fe8),
	.w7(32'hbc0ba2b5),
	.w8(32'h3c884132),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce6218a),
	.w1(32'hbb42dcb5),
	.w2(32'hbd53820f),
	.w3(32'h3ca86950),
	.w4(32'h3b4fe076),
	.w5(32'hbca3a1a7),
	.w6(32'hbc672e28),
	.w7(32'hbd1af382),
	.w8(32'hbac68ae2),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd31fb4),
	.w1(32'h3a9f6bc3),
	.w2(32'h3b218bde),
	.w3(32'hbb0cdf9c),
	.w4(32'h39b94561),
	.w5(32'h399e34f7),
	.w6(32'h3b124dd2),
	.w7(32'h3a3fec1f),
	.w8(32'hbca9af05),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd6a8325),
	.w1(32'hbc10261e),
	.w2(32'h3d352ae8),
	.w3(32'hbd18b769),
	.w4(32'hbc2400f9),
	.w5(32'h3c93e86b),
	.w6(32'h3b1b261f),
	.w7(32'h3cd3cfe3),
	.w8(32'h3cbd23bf),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d1faa5f),
	.w1(32'hbab51dab),
	.w2(32'hbd38cf0c),
	.w3(32'h3d0660a2),
	.w4(32'h3bff6346),
	.w5(32'hbcd15f97),
	.w6(32'hbc0ed430),
	.w7(32'hbd251b5a),
	.w8(32'h3bf64bb9),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca52131),
	.w1(32'h3b2431a5),
	.w2(32'hbc18d8b7),
	.w3(32'h3c3c4423),
	.w4(32'h3b28a234),
	.w5(32'hbb7977f0),
	.w6(32'hbb23231f),
	.w7(32'hbbadbd97),
	.w8(32'hb990e696),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f28f60),
	.w1(32'hba35f804),
	.w2(32'hbab28e0b),
	.w3(32'hbab5d985),
	.w4(32'hbac80550),
	.w5(32'hbac927aa),
	.w6(32'hbaaa874f),
	.w7(32'hba3d3d2b),
	.w8(32'hbb387151),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6bf480),
	.w1(32'hba6bb9bd),
	.w2(32'hb948051a),
	.w3(32'hbb69537f),
	.w4(32'hb9318727),
	.w5(32'hbae443b3),
	.w6(32'h3aa090ae),
	.w7(32'hba3d4302),
	.w8(32'hb9875d7c),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb861c3df),
	.w1(32'h392741f7),
	.w2(32'h39a4b152),
	.w3(32'h39c2d9a3),
	.w4(32'h3a2fe6e4),
	.w5(32'h39c01127),
	.w6(32'hb9bd106c),
	.w7(32'h37e28cea),
	.w8(32'h3a17f13d),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d34225),
	.w1(32'hb56ffcb4),
	.w2(32'h38f7a5bc),
	.w3(32'h39b3c240),
	.w4(32'h37c6b97a),
	.w5(32'h38a7a8b3),
	.w6(32'hb9925480),
	.w7(32'h38236b6c),
	.w8(32'h3915d50e),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f0c2f6),
	.w1(32'hb9c45234),
	.w2(32'hb849da86),
	.w3(32'h3a7bf6c9),
	.w4(32'h396d6db8),
	.w5(32'h3a78efcb),
	.w6(32'hba2c19de),
	.w7(32'hb99b2dcb),
	.w8(32'hbac93c32),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb40b3da),
	.w1(32'hbb4a72d1),
	.w2(32'hbbada6df),
	.w3(32'hbac86347),
	.w4(32'h3963f4e0),
	.w5(32'hb9e30887),
	.w6(32'hbb1a66d1),
	.w7(32'hbabb7a2d),
	.w8(32'h39b824cc),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d8cff6),
	.w1(32'hba5fa70d),
	.w2(32'hb6c9f55d),
	.w3(32'hb9157eba),
	.w4(32'hb98f92ed),
	.w5(32'h3981d214),
	.w6(32'hbaa5920e),
	.w7(32'h399cef84),
	.w8(32'h399dfef5),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d602ca),
	.w1(32'hb984d887),
	.w2(32'h399b5073),
	.w3(32'hba5aaf7f),
	.w4(32'hb98d835f),
	.w5(32'h39b2d03c),
	.w6(32'h39e4a5f0),
	.w7(32'h3ac13b42),
	.w8(32'h39b8f394),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a57f537),
	.w1(32'h37a74e9b),
	.w2(32'h39eed521),
	.w3(32'h3a5ef58f),
	.w4(32'h39b7f299),
	.w5(32'h3a30fcef),
	.w6(32'hb95fd033),
	.w7(32'h39629b96),
	.w8(32'hb953d938),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3941b90a),
	.w1(32'hb94d969a),
	.w2(32'h38f25ee3),
	.w3(32'h389f2c2d),
	.w4(32'hb9860369),
	.w5(32'hb9725b52),
	.w6(32'hb9eb0670),
	.w7(32'hb9c9d079),
	.w8(32'hba17f351),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb84dabb7),
	.w1(32'hba064ef7),
	.w2(32'hb95c3839),
	.w3(32'hb8ddd103),
	.w4(32'hb9ed009b),
	.w5(32'hb9b718f5),
	.w6(32'hba890730),
	.w7(32'hba5f7b4c),
	.w8(32'hba1655dc),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6b0480),
	.w1(32'hbb295e92),
	.w2(32'hbb5f7375),
	.w3(32'hba434f17),
	.w4(32'hbad51e68),
	.w5(32'hbabe5e1e),
	.w6(32'hb99c4653),
	.w7(32'hb9cc3b0b),
	.w8(32'hb9676980),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7b58ad),
	.w1(32'hba4db0c5),
	.w2(32'hba69557b),
	.w3(32'hba56e5ea),
	.w4(32'hba14c123),
	.w5(32'hba07930a),
	.w6(32'hba600084),
	.w7(32'hb9110cd7),
	.w8(32'h39a1b453),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad504ad),
	.w1(32'hbb016d41),
	.w2(32'hbb5d169d),
	.w3(32'hba0d275c),
	.w4(32'hb967ecb8),
	.w5(32'hbaf4c684),
	.w6(32'hba2b9f7b),
	.w7(32'hbb1f05c8),
	.w8(32'hbab47319),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeee102),
	.w1(32'hbb674b32),
	.w2(32'hbb1e085d),
	.w3(32'hbac304a5),
	.w4(32'hbb5b7082),
	.w5(32'hbb01d088),
	.w6(32'hbb05c1b0),
	.w7(32'hba92b7b6),
	.w8(32'hb9fb8644),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb124d97),
	.w1(32'hbac1f2c1),
	.w2(32'hb99cb5a1),
	.w3(32'h39c530c5),
	.w4(32'h37af3e3c),
	.w5(32'h3a33a229),
	.w6(32'hba3a5d93),
	.w7(32'hba9181f9),
	.w8(32'hba9c78c6),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6c5eac),
	.w1(32'hbb0d8e9e),
	.w2(32'hbb1b3123),
	.w3(32'hb9f2ccb5),
	.w4(32'hbafd7103),
	.w5(32'hbac25a65),
	.w6(32'h3a33b245),
	.w7(32'hb9713a6c),
	.w8(32'h3a8890df),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3946ea79),
	.w1(32'h378c40eb),
	.w2(32'h3a81b438),
	.w3(32'h3981edff),
	.w4(32'h393de942),
	.w5(32'h3a732fd4),
	.w6(32'h3aa619be),
	.w7(32'h3b068579),
	.w8(32'hba965d17),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0d52e7),
	.w1(32'hba3f04c8),
	.w2(32'hbaa04109),
	.w3(32'hba498d31),
	.w4(32'hba99debf),
	.w5(32'hba4d69df),
	.w6(32'hba349155),
	.w7(32'hba91a01e),
	.w8(32'h3a45e9e6),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4013fd),
	.w1(32'hbb241cb3),
	.w2(32'hbade6140),
	.w3(32'h39b0fc34),
	.w4(32'h392e3211),
	.w5(32'hb9c84b90),
	.w6(32'hba90d9ba),
	.w7(32'hbb28cc19),
	.w8(32'h3a408591),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e66809),
	.w1(32'hba10dd5a),
	.w2(32'hba18936d),
	.w3(32'h3a7b38ce),
	.w4(32'h39642413),
	.w5(32'h3a3a839c),
	.w6(32'hba68a1a0),
	.w7(32'hb9db79e5),
	.w8(32'h3a0a77a3),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8d3b57),
	.w1(32'h3999ca73),
	.w2(32'h39ec653a),
	.w3(32'h3a95d47a),
	.w4(32'h3a3bad38),
	.w5(32'h3a1e738a),
	.w6(32'h398292bc),
	.w7(32'h39f571d5),
	.w8(32'hb80dbb88),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf2b089),
	.w1(32'hbafd5f5a),
	.w2(32'hba969a53),
	.w3(32'hb95fa596),
	.w4(32'hbb1ad917),
	.w5(32'hbafbdeaa),
	.w6(32'h3a87a9f8),
	.w7(32'h3ae1a29a),
	.w8(32'hb968f484),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule