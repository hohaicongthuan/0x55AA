module layer_8_featuremap_16(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c497c6a),
	.w1(32'hbbbf5404),
	.w2(32'hbb3f808c),
	.w3(32'hbc1fb2f8),
	.w4(32'hbca08337),
	.w5(32'h3bd71db9),
	.w6(32'hbc05ed92),
	.w7(32'hbac474fd),
	.w8(32'h3c4b7f28),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8d3c474),
	.w1(32'hbbeca092),
	.w2(32'h3bf0a6ae),
	.w3(32'h3c1ade2d),
	.w4(32'h3c4b9e71),
	.w5(32'h3b0c4e78),
	.w6(32'h3be8de6a),
	.w7(32'hbb7420c5),
	.w8(32'h3c554f1a),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ca0e413),
	.w1(32'hbc600099),
	.w2(32'hb847480b),
	.w3(32'hbc554f27),
	.w4(32'h3a245fd2),
	.w5(32'hbb4d9a8e),
	.w6(32'h3c82c703),
	.w7(32'h3c66448e),
	.w8(32'h3ab744a6),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acc14ba),
	.w1(32'h3c8a6413),
	.w2(32'h3b83e5c7),
	.w3(32'h3be25de4),
	.w4(32'h3b42cbbb),
	.w5(32'h3c6f5776),
	.w6(32'hbbad9c2f),
	.w7(32'h3b9fab61),
	.w8(32'h3c3df84f),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c13cf36),
	.w1(32'hbb268e7b),
	.w2(32'h3a414a3a),
	.w3(32'h3bb81d99),
	.w4(32'h3bb21c6f),
	.w5(32'h3a5f010b),
	.w6(32'h3a09a688),
	.w7(32'hbbc910e6),
	.w8(32'h3b2efbed),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfb4633),
	.w1(32'hbcc379d3),
	.w2(32'hbc0d9be9),
	.w3(32'h3cb4ec2c),
	.w4(32'h3b8a828e),
	.w5(32'h38f1ff3e),
	.w6(32'h3c43a7e5),
	.w7(32'hbc0d27d1),
	.w8(32'h3b7eb230),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb20b79e),
	.w1(32'hbc300ee2),
	.w2(32'h3b3c562d),
	.w3(32'h3d0fb473),
	.w4(32'hbace930e),
	.w5(32'h3a7da69f),
	.w6(32'h3ad5ddd9),
	.w7(32'h3c72b509),
	.w8(32'h3af6b489),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba98eab2),
	.w1(32'h3c0d83d7),
	.w2(32'h3bb94881),
	.w3(32'h3bfe49e6),
	.w4(32'hbbcf6fe4),
	.w5(32'h3c8c7c3a),
	.w6(32'hbb9c9f4d),
	.w7(32'h3c914749),
	.w8(32'hbbda1807),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8b5671),
	.w1(32'hbb04d758),
	.w2(32'hbb434afc),
	.w3(32'h3c80c32f),
	.w4(32'hbb99afe8),
	.w5(32'h3b3c35d4),
	.w6(32'hbac2006e),
	.w7(32'hbc9933c5),
	.w8(32'hbc565c80),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f06055),
	.w1(32'hbad34673),
	.w2(32'hbbbb0dea),
	.w3(32'h3ae87d5d),
	.w4(32'hbc38c8ba),
	.w5(32'hbbe27daa),
	.w6(32'hbbb2fa78),
	.w7(32'hbc845fae),
	.w8(32'h3b9cdc4b),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcd91b3),
	.w1(32'h3ca3976b),
	.w2(32'hbc34cd09),
	.w3(32'hba8d1ef5),
	.w4(32'hbc188553),
	.w5(32'h3b814346),
	.w6(32'h3b6dd1e5),
	.w7(32'hbc2f52ea),
	.w8(32'hbcb0252e),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb10c87c),
	.w1(32'h3c63212e),
	.w2(32'h3a98699f),
	.w3(32'h3b5f3a58),
	.w4(32'hbc4bf6d4),
	.w5(32'hbc3305e8),
	.w6(32'hbbeea66e),
	.w7(32'h3cddf37e),
	.w8(32'h3bb7a0e3),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d76a1e),
	.w1(32'h3bef3a0a),
	.w2(32'hbc104aef),
	.w3(32'hbc91fea3),
	.w4(32'hbaa81a7a),
	.w5(32'h39a415fc),
	.w6(32'h3c8e37d5),
	.w7(32'h3c0e00e1),
	.w8(32'hbc1246cb),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc438d6e),
	.w1(32'h3b4b78a5),
	.w2(32'hbcb4cc88),
	.w3(32'h3b1f7848),
	.w4(32'hbbb770d2),
	.w5(32'hbbabf98b),
	.w6(32'hbb8758ca),
	.w7(32'h3cd1fb47),
	.w8(32'h3b7bfea9),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba61dc16),
	.w1(32'hbbcf68c6),
	.w2(32'hbcf8813c),
	.w3(32'hbbb25f68),
	.w4(32'hbb9b5b95),
	.w5(32'h3c5f54fc),
	.w6(32'h3d09cfab),
	.w7(32'hbc388eb8),
	.w8(32'h3bf825a9),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb97e8e),
	.w1(32'h3b9cda63),
	.w2(32'h3ba18a26),
	.w3(32'hbc25f019),
	.w4(32'hbb7fe0b0),
	.w5(32'hbc2a3fdc),
	.w6(32'h39bb4907),
	.w7(32'hb99ede46),
	.w8(32'hbb18b046),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf88ea7),
	.w1(32'h3b85c3ef),
	.w2(32'h3a368658),
	.w3(32'h3b01b55c),
	.w4(32'hbbfcc74f),
	.w5(32'h3cc5dbf3),
	.w6(32'hbc4f3a43),
	.w7(32'hba49f47f),
	.w8(32'hbb4b1674),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2e3c4b),
	.w1(32'h3b678385),
	.w2(32'hbc847e0d),
	.w3(32'h3b3ebde1),
	.w4(32'hbc3b53ef),
	.w5(32'hbb9eefde),
	.w6(32'hbc4dff78),
	.w7(32'h3b42b97c),
	.w8(32'hb7c73a62),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0fa363),
	.w1(32'hbb2f4599),
	.w2(32'hbc312dac),
	.w3(32'hbbc230eb),
	.w4(32'hbb7fa78e),
	.w5(32'hbbfa0bbf),
	.w6(32'h3aa23509),
	.w7(32'h3af16a28),
	.w8(32'hbbe2354b),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cb71b9),
	.w1(32'hbccfba96),
	.w2(32'h3bd6b27c),
	.w3(32'h3b950110),
	.w4(32'h3c887a5c),
	.w5(32'hbb15c92c),
	.w6(32'hb9fca74e),
	.w7(32'hbaf5b7a2),
	.w8(32'h3c3cd1f8),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb717e4d8),
	.w1(32'hbcca86d7),
	.w2(32'hbc1a784c),
	.w3(32'hbc213305),
	.w4(32'h3bcf1f46),
	.w5(32'h3ba54dad),
	.w6(32'hbb588431),
	.w7(32'hbb432c80),
	.w8(32'h3b29f8d8),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbd1fb342),
	.w1(32'h3c646036),
	.w2(32'hbb26c243),
	.w3(32'h3bb01d02),
	.w4(32'hbc0c9bf8),
	.w5(32'hbc0a2e5e),
	.w6(32'h3ba0e44e),
	.w7(32'hbc6b1178),
	.w8(32'h3c0f1956),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc60fb3b),
	.w1(32'hbb8766dd),
	.w2(32'hbb5fbef7),
	.w3(32'hbbd4b076),
	.w4(32'hba1c5372),
	.w5(32'hbb0de6b0),
	.w6(32'hbb124786),
	.w7(32'hbc48be1f),
	.w8(32'h3a86b0fd),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbc7840),
	.w1(32'hbc1af731),
	.w2(32'hbca05ee2),
	.w3(32'hbcd08723),
	.w4(32'hbc9a97e5),
	.w5(32'hbbc786a6),
	.w6(32'h39e02017),
	.w7(32'hbc0d549f),
	.w8(32'h3b94ea3c),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc61fd9),
	.w1(32'h3b17f546),
	.w2(32'hb8c04e08),
	.w3(32'hbb14a808),
	.w4(32'h3c69a856),
	.w5(32'hbc9411d8),
	.w6(32'h39f96af1),
	.w7(32'h3c3a4f93),
	.w8(32'hbb2c2463),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b854a44),
	.w1(32'h3b786066),
	.w2(32'h3b994cbf),
	.w3(32'h3c4e895c),
	.w4(32'hbc878462),
	.w5(32'h3aa5b96b),
	.w6(32'hbab97e68),
	.w7(32'hbc3eb379),
	.w8(32'h398cf406),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbceb1d6),
	.w1(32'h3c1f87da),
	.w2(32'hbbb24daa),
	.w3(32'hbb66838d),
	.w4(32'hbcb129c8),
	.w5(32'hbc570dc2),
	.w6(32'hbb8bbcd9),
	.w7(32'hbb20b49b),
	.w8(32'h3bb1f947),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b139949),
	.w1(32'hbb7e1c24),
	.w2(32'h3c159cad),
	.w3(32'h3c98d3be),
	.w4(32'hbc59c098),
	.w5(32'hbabc9057),
	.w6(32'hbc4c0b93),
	.w7(32'hbc6584f5),
	.w8(32'hbceb0ef8),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8e67e3),
	.w1(32'h3d2032f6),
	.w2(32'hbb818a28),
	.w3(32'hbc2b0f5f),
	.w4(32'h37a52da3),
	.w5(32'h3c482a0e),
	.w6(32'hbb0e4ab1),
	.w7(32'hbc80eb6c),
	.w8(32'h3cf8e3a8),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb45f83a),
	.w1(32'hbc6aa3e1),
	.w2(32'h3cc909d6),
	.w3(32'hbc77c983),
	.w4(32'hbc7be98b),
	.w5(32'hbc40130b),
	.w6(32'hbca65093),
	.w7(32'hb9383ef2),
	.w8(32'h3c635084),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba2f2d3),
	.w1(32'h3cef81fb),
	.w2(32'hbc4890ca),
	.w3(32'hbbb668e0),
	.w4(32'hbc492c19),
	.w5(32'hbd45d6ef),
	.w6(32'hbca8fe84),
	.w7(32'h3c70719a),
	.w8(32'h3a93cf15),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0c65b4),
	.w1(32'h3c2f50ae),
	.w2(32'h3b8474ca),
	.w3(32'hbd0cb2a1),
	.w4(32'hbcbb8f7c),
	.w5(32'hbc714650),
	.w6(32'hbc825123),
	.w7(32'h3b6a6d4f),
	.w8(32'hbb22218d),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc190ebd),
	.w1(32'h3d576714),
	.w2(32'h3addb27c),
	.w3(32'hbd1099df),
	.w4(32'hbc320de5),
	.w5(32'hbc88371c),
	.w6(32'hbcd1a2eb),
	.w7(32'h3b370528),
	.w8(32'h3aa06dbd),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c169ed7),
	.w1(32'h3c591fb1),
	.w2(32'h3c9dc570),
	.w3(32'hbbe587fc),
	.w4(32'hbb5df2ca),
	.w5(32'hbabd04d3),
	.w6(32'h3aa79ce2),
	.w7(32'hbb6c9585),
	.w8(32'h39abe033),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bee774c),
	.w1(32'hbcd3cde7),
	.w2(32'hbc401521),
	.w3(32'hbc6fe7b7),
	.w4(32'h3cef2d70),
	.w5(32'h3c880117),
	.w6(32'hbc3bb76d),
	.w7(32'hbca687cb),
	.w8(32'hbc93d5f9),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc6531f),
	.w1(32'hbb9738dd),
	.w2(32'hbb2da829),
	.w3(32'h39ee01c6),
	.w4(32'h3b79c866),
	.w5(32'h3c931244),
	.w6(32'hbb9a8fc0),
	.w7(32'hbaad47da),
	.w8(32'h3c82e186),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca2c041),
	.w1(32'hbc940d71),
	.w2(32'hbaa3306c),
	.w3(32'hbc30b81b),
	.w4(32'hbac48adb),
	.w5(32'h38678c72),
	.w6(32'h3c1c83ae),
	.w7(32'h3cba78d7),
	.w8(32'hbc5fbc5a),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c08bc8d),
	.w1(32'hb95f756a),
	.w2(32'hbd07ae75),
	.w3(32'hba8a26ed),
	.w4(32'hb888dc3e),
	.w5(32'hbd19b9f2),
	.w6(32'hba9c93e1),
	.w7(32'hbca792f7),
	.w8(32'h3cfeaceb),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf7c20a),
	.w1(32'hbc493221),
	.w2(32'hbaca873d),
	.w3(32'hbc479c3c),
	.w4(32'hbc54fd44),
	.w5(32'h3c4b7d53),
	.w6(32'h3c50c754),
	.w7(32'hbbdb446f),
	.w8(32'hbc5c9b5e),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2bc62b),
	.w1(32'h3ba09977),
	.w2(32'hba11b09e),
	.w3(32'h3cbf6c68),
	.w4(32'h3d3de383),
	.w5(32'hbc8c559a),
	.w6(32'hbb159300),
	.w7(32'hbc33f6c8),
	.w8(32'h3c4d116d),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d2f5c46),
	.w1(32'h3d3d4147),
	.w2(32'h3bc04225),
	.w3(32'hba5f4e57),
	.w4(32'h399412c6),
	.w5(32'hbd26244d),
	.w6(32'h3c13645e),
	.w7(32'hbc024868),
	.w8(32'h3b157163),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb808ecd),
	.w1(32'hbb6f1142),
	.w2(32'hbb917cda),
	.w3(32'hba400d32),
	.w4(32'hb8ab44d6),
	.w5(32'hba0eaa7e),
	.w6(32'h3bc42db2),
	.w7(32'hbb29bad1),
	.w8(32'hb9f12519),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c442166),
	.w1(32'hb9987d5d),
	.w2(32'h3c427a63),
	.w3(32'hbb367c2c),
	.w4(32'h3c01f892),
	.w5(32'h3b1c839d),
	.w6(32'h3bbd036f),
	.w7(32'hbb2ab044),
	.w8(32'hb925d6d8),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2cdee3),
	.w1(32'hbbbe260f),
	.w2(32'h3a898f04),
	.w3(32'h3b1f05e5),
	.w4(32'hbb6b0fa8),
	.w5(32'h3a121fa9),
	.w6(32'hbb2d9c69),
	.w7(32'hbb901555),
	.w8(32'hbba23010),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a452453),
	.w1(32'h3b967d3f),
	.w2(32'h3b425fd7),
	.w3(32'hbba3f917),
	.w4(32'hbac495b3),
	.w5(32'hbb60b258),
	.w6(32'hbbb00a12),
	.w7(32'h3b98821f),
	.w8(32'hbb1c3bdf),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcdd1cb),
	.w1(32'h3b0079c3),
	.w2(32'h39c357ae),
	.w3(32'h39ba5a40),
	.w4(32'hbb627ed2),
	.w5(32'hb7ce1202),
	.w6(32'h3b792387),
	.w7(32'hb9ca0ce3),
	.w8(32'h3a29695d),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c04ec10),
	.w1(32'h3ac5d25d),
	.w2(32'hba839f35),
	.w3(32'hbb035777),
	.w4(32'hbbbf1f18),
	.w5(32'h3a32a869),
	.w6(32'h3bf43e73),
	.w7(32'hbb883ca0),
	.w8(32'h3bc0ebf4),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb100d41),
	.w1(32'hbb8a7c36),
	.w2(32'hbabd1ece),
	.w3(32'h3c746a3f),
	.w4(32'h3b070a5e),
	.w5(32'h3b8b6988),
	.w6(32'hbb6dec90),
	.w7(32'h3a84829a),
	.w8(32'h3b229caa),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b6b82),
	.w1(32'h3a841778),
	.w2(32'hbb58dfe1),
	.w3(32'h3b57dde1),
	.w4(32'h3bbbfdce),
	.w5(32'h3adac312),
	.w6(32'h3c088467),
	.w7(32'hbb8062f5),
	.w8(32'h3c1779d9),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbffd89e),
	.w1(32'h3ad7e892),
	.w2(32'h3b38f5d8),
	.w3(32'hbbac27d4),
	.w4(32'hbb47f62c),
	.w5(32'h3c2fe271),
	.w6(32'h3c7916aa),
	.w7(32'h39d18c98),
	.w8(32'hbbb98e7b),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbe98e8),
	.w1(32'h3c18fc0b),
	.w2(32'h3a6a6e5f),
	.w3(32'hb91d8466),
	.w4(32'hb9f6332f),
	.w5(32'hbaf1525c),
	.w6(32'h3ba4fe1f),
	.w7(32'h3b2b0f53),
	.w8(32'h3a8976bc),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadb2f26),
	.w1(32'hba542eec),
	.w2(32'h38d5e9f3),
	.w3(32'hbbb44743),
	.w4(32'hbb1efc70),
	.w5(32'hb9ae4137),
	.w6(32'hbb80ed50),
	.w7(32'h3b591e53),
	.w8(32'hba7c197c),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb005f99),
	.w1(32'h3b500d66),
	.w2(32'hbb1d67c5),
	.w3(32'h3ba23e6e),
	.w4(32'hbbbabbcd),
	.w5(32'h3c8a08b0),
	.w6(32'hba9feb36),
	.w7(32'h3a87df1f),
	.w8(32'h3c3f8680),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcce89b),
	.w1(32'hbb4a0583),
	.w2(32'hba66847c),
	.w3(32'hbbfeffe4),
	.w4(32'h3a6b77f4),
	.w5(32'hb91dceb9),
	.w6(32'hbbb01729),
	.w7(32'hbaa17973),
	.w8(32'h3a9c3231),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6ad93e),
	.w1(32'h39c49e68),
	.w2(32'hbb1f68d2),
	.w3(32'h3a831d15),
	.w4(32'hbbac0991),
	.w5(32'h3a812f4d),
	.w6(32'h38912a0d),
	.w7(32'h3bf91fab),
	.w8(32'hba5942e6),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1d9956),
	.w1(32'hbae21a4c),
	.w2(32'hbaa43d37),
	.w3(32'hbb2ebb4e),
	.w4(32'h3bb6496f),
	.w5(32'h3beaf446),
	.w6(32'h3b246920),
	.w7(32'hbb0143c5),
	.w8(32'hbb8d58d9),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93712f0),
	.w1(32'hb8d1b0ab),
	.w2(32'h3b29c500),
	.w3(32'hb98ef1de),
	.w4(32'h3aea4b66),
	.w5(32'h3835452f),
	.w6(32'h3c9c8361),
	.w7(32'h3a0fff21),
	.w8(32'h3b4f679b),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3891d1f0),
	.w1(32'h3a10731e),
	.w2(32'h394c3500),
	.w3(32'hba45141e),
	.w4(32'hba9ef656),
	.w5(32'h38d33d4f),
	.w6(32'hbad4e651),
	.w7(32'hba504fda),
	.w8(32'h3b1a389c),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb902d528),
	.w1(32'h3a8438a2),
	.w2(32'hbb1dc579),
	.w3(32'hb9b17694),
	.w4(32'hbbd2fc6b),
	.w5(32'hbb657da7),
	.w6(32'h3888144b),
	.w7(32'h3ac4eb64),
	.w8(32'h3ae3c4aa),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d276f9),
	.w1(32'h39afc1d5),
	.w2(32'hbb463c78),
	.w3(32'hb6210256),
	.w4(32'h3a175712),
	.w5(32'hbb2568ed),
	.w6(32'h3b4390d1),
	.w7(32'hb7a09dfb),
	.w8(32'hbb898587),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaac2f4),
	.w1(32'hbb9ec86e),
	.w2(32'h3b15ed34),
	.w3(32'hba6e7ff7),
	.w4(32'h3b4950e5),
	.w5(32'hbb0dbee4),
	.w6(32'hba55e869),
	.w7(32'hb9e26e49),
	.w8(32'hbb3670c2),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a4805b),
	.w1(32'h38e12567),
	.w2(32'h3a92b92b),
	.w3(32'h3aa85b05),
	.w4(32'hbad5667d),
	.w5(32'h3a4671cf),
	.w6(32'h3a30d22b),
	.w7(32'hba1f14eb),
	.w8(32'h3a1712ba),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b88d8d8),
	.w1(32'h3a1a079a),
	.w2(32'h3ae2cad3),
	.w3(32'h3bb05027),
	.w4(32'hba5ca80b),
	.w5(32'h3ad6a768),
	.w6(32'hbbdca4b9),
	.w7(32'h3ac98145),
	.w8(32'h3a7c7919),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba09b275),
	.w1(32'h3a09654d),
	.w2(32'h3b072374),
	.w3(32'h3be83af6),
	.w4(32'h3b3a5956),
	.w5(32'h3969c535),
	.w6(32'hb938e7c1),
	.w7(32'h3b263e75),
	.w8(32'h3af9bc60),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c074d1e),
	.w1(32'h3a926171),
	.w2(32'h3adf455e),
	.w3(32'h39fd7880),
	.w4(32'h3b3983b8),
	.w5(32'hba591842),
	.w6(32'hbb45b40c),
	.w7(32'h39c0372e),
	.w8(32'h39bc5fd8),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbc095b),
	.w1(32'hba268311),
	.w2(32'hbb6e4338),
	.w3(32'hb976b58a),
	.w4(32'h3a4fd546),
	.w5(32'h3a8abf4c),
	.w6(32'hbb3865bd),
	.w7(32'hbb4b7d0d),
	.w8(32'h38b936d1),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9265ef),
	.w1(32'h395e5756),
	.w2(32'h3b71134c),
	.w3(32'hb814e1e6),
	.w4(32'h3b15c262),
	.w5(32'h3a15eec3),
	.w6(32'h3a08d780),
	.w7(32'hbb9c9d13),
	.w8(32'h3b472f4c),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbfc122),
	.w1(32'hbab9973b),
	.w2(32'h3a4dacff),
	.w3(32'h3b9cd14f),
	.w4(32'hbb8d6bb3),
	.w5(32'h3bedcadf),
	.w6(32'h3b499c84),
	.w7(32'h3a5b00dd),
	.w8(32'hb99bce1e),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba69b1fa),
	.w1(32'hbb032e30),
	.w2(32'hb9957bd6),
	.w3(32'hba101a1f),
	.w4(32'hbac24969),
	.w5(32'hba20c8da),
	.w6(32'h3be491c1),
	.w7(32'h3a2fea2e),
	.w8(32'hbb7afbed),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5913f1),
	.w1(32'hbad0742b),
	.w2(32'h3a907112),
	.w3(32'hbb0da513),
	.w4(32'h3b3f67db),
	.w5(32'hba40551d),
	.w6(32'hbb22ccab),
	.w7(32'hbae4e8a1),
	.w8(32'hbb5ea985),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b74c7db),
	.w1(32'h3a9dc0d7),
	.w2(32'h3aca338a),
	.w3(32'h3accc0b9),
	.w4(32'h3c548dac),
	.w5(32'h3aba6949),
	.w6(32'h3b187df3),
	.w7(32'hbb7d96c0),
	.w8(32'h3baad571),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b8f0ba),
	.w1(32'hba4080ab),
	.w2(32'h3ba650da),
	.w3(32'h3ba6cfaf),
	.w4(32'hba1c2742),
	.w5(32'h3a070c9a),
	.w6(32'hbac09f4b),
	.w7(32'h3ab0618e),
	.w8(32'hba7052ad),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7f94c5),
	.w1(32'h3a091d40),
	.w2(32'hbbcf0a50),
	.w3(32'h3a92ad53),
	.w4(32'h36062f85),
	.w5(32'h396bcf30),
	.w6(32'h3a40a45e),
	.w7(32'hba8ba058),
	.w8(32'hbb14d145),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4d0c8d),
	.w1(32'hba9501bd),
	.w2(32'hbb46b0f8),
	.w3(32'hbbb84af8),
	.w4(32'h3afcfbb6),
	.w5(32'hba555e24),
	.w6(32'hbb409a7b),
	.w7(32'hba63e52b),
	.w8(32'h3ac2ffd8),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad1f0de),
	.w1(32'hbb2d8f74),
	.w2(32'h3bd59c7e),
	.w3(32'hbbb2b1c6),
	.w4(32'h3b7d8f3c),
	.w5(32'h3ae9a0d5),
	.w6(32'h3970f8ca),
	.w7(32'hb98f87d1),
	.w8(32'hba62be94),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba18c682),
	.w1(32'hbb5d06c8),
	.w2(32'hba1c576f),
	.w3(32'hbac787f7),
	.w4(32'hbaeb894f),
	.w5(32'hbaad2e83),
	.w6(32'h3a28a83d),
	.w7(32'hbb3590be),
	.w8(32'h3a258ec0),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b29643c),
	.w1(32'h3bc6c6d9),
	.w2(32'hbb460923),
	.w3(32'hbb192c48),
	.w4(32'hbbc22940),
	.w5(32'h3ad4f5e2),
	.w6(32'h39986581),
	.w7(32'h3ac3a62b),
	.w8(32'h391cd6e2),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b24de2d),
	.w1(32'h3baac40d),
	.w2(32'h3a08f3df),
	.w3(32'h3a6f4caf),
	.w4(32'hba1fcbf6),
	.w5(32'h3a83b41c),
	.w6(32'hbb61f363),
	.w7(32'h3b139cb4),
	.w8(32'hbbd7f8ac),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8a97e7a),
	.w1(32'hb9be36a9),
	.w2(32'hba949c90),
	.w3(32'h3b81612a),
	.w4(32'hbba997a1),
	.w5(32'hb98059cf),
	.w6(32'h3bc70111),
	.w7(32'hbb21044d),
	.w8(32'h3a18e3a4),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e56485),
	.w1(32'h39331dd4),
	.w2(32'h3a0c9e71),
	.w3(32'hb881912c),
	.w4(32'h37aa4f55),
	.w5(32'hbb47e31c),
	.w6(32'hbb9fe311),
	.w7(32'hbb3d3c5a),
	.w8(32'hbabf0870),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb6fb3f08),
	.w1(32'hbb634cb3),
	.w2(32'h388bf309),
	.w3(32'h39e7f2d9),
	.w4(32'hbac580dc),
	.w5(32'hbbbd3cbb),
	.w6(32'h39abfd3d),
	.w7(32'h3b338e28),
	.w8(32'h3b079d69),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a92c6b6),
	.w1(32'h3bde8e0b),
	.w2(32'hbb618025),
	.w3(32'hb877059d),
	.w4(32'h3b913822),
	.w5(32'h3a085414),
	.w6(32'hbb4d711a),
	.w7(32'hba9e685c),
	.w8(32'h3aa47e5d),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc315ca0),
	.w1(32'hbadd2c9a),
	.w2(32'h3ab80127),
	.w3(32'hba0dafbd),
	.w4(32'hba8dffc1),
	.w5(32'h3a1490a9),
	.w6(32'hb84a3564),
	.w7(32'hbbd0f531),
	.w8(32'hb9eeb41b),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b799e65),
	.w1(32'hbb557a8f),
	.w2(32'hbabdb9f3),
	.w3(32'hbb2593bc),
	.w4(32'hba386fc7),
	.w5(32'h3c9c5489),
	.w6(32'hbbe21534),
	.w7(32'h3a929ff6),
	.w8(32'hbad581a6),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9c3016),
	.w1(32'h3bbcbbf9),
	.w2(32'h3b13ad04),
	.w3(32'h3b32bb32),
	.w4(32'hbba3c62d),
	.w5(32'h3c132dd5),
	.w6(32'h38bc8f04),
	.w7(32'h39b30a0e),
	.w8(32'hbc8c8629),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7b5932e),
	.w1(32'hba60ff2b),
	.w2(32'h3be10f98),
	.w3(32'hbbf74955),
	.w4(32'hbb5a24a3),
	.w5(32'hbd035c8a),
	.w6(32'hbb14eee5),
	.w7(32'hb78a9240),
	.w8(32'hbb2b5e88),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb216ed4),
	.w1(32'hb98cba72),
	.w2(32'hbbab9759),
	.w3(32'hbbdc9486),
	.w4(32'hbaabad34),
	.w5(32'hbcaabfa5),
	.w6(32'hbc4ffc64),
	.w7(32'h3b125bf1),
	.w8(32'h3aa1e9af),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8f80a4),
	.w1(32'h3bd19d01),
	.w2(32'h3b822c92),
	.w3(32'h3c85314c),
	.w4(32'hbc376789),
	.w5(32'hb9293b7f),
	.w6(32'h3a3b4fc0),
	.w7(32'h37a73b4f),
	.w8(32'h3a94b20a),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba0f5ed),
	.w1(32'h3bd4fe9e),
	.w2(32'hbac3b30b),
	.w3(32'h3bbad86f),
	.w4(32'hba054673),
	.w5(32'h3b41350f),
	.w6(32'h3799fcfc),
	.w7(32'h3b8e4c73),
	.w8(32'hbc50760c),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb973b76),
	.w1(32'h3bd73bd2),
	.w2(32'hba933a82),
	.w3(32'h3b846305),
	.w4(32'h3a162dd0),
	.w5(32'hbc191a7b),
	.w6(32'h3abd20a2),
	.w7(32'h3b908e69),
	.w8(32'h3b0982a1),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc501d59),
	.w1(32'hbbe615f0),
	.w2(32'hbc3e4fb7),
	.w3(32'hba911686),
	.w4(32'h3bc4d56a),
	.w5(32'hbb448c44),
	.w6(32'hbb2b78a6),
	.w7(32'hbc2dd1f9),
	.w8(32'h39477dd2),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8c492a),
	.w1(32'hbc1084d0),
	.w2(32'h3cbc125d),
	.w3(32'h3b0ab20a),
	.w4(32'h3c67a2a0),
	.w5(32'h3cea908c),
	.w6(32'h3b73bed7),
	.w7(32'hba5bf8b9),
	.w8(32'h3b850ce8),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4d0a58),
	.w1(32'hbb9aedf1),
	.w2(32'h3bfcb845),
	.w3(32'hbbda0e21),
	.w4(32'h3bc5d5b8),
	.w5(32'hbc38069a),
	.w6(32'hb9bfadda),
	.w7(32'hbb40c0bf),
	.w8(32'hbbcc5844),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbdbe78),
	.w1(32'hb9b6beed),
	.w2(32'h3c609ca1),
	.w3(32'h3c8d0f03),
	.w4(32'hbbc9bf83),
	.w5(32'h3c940620),
	.w6(32'hbb285b88),
	.w7(32'hb9960e75),
	.w8(32'hbc1c752c),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b76e9a6),
	.w1(32'h392ea552),
	.w2(32'h3c886fb3),
	.w3(32'hb6635ae2),
	.w4(32'hbc563e54),
	.w5(32'hbc52de27),
	.w6(32'hbc98aaaf),
	.w7(32'h3add04c1),
	.w8(32'hbc2d354b),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3caec64c),
	.w1(32'h3b038ceb),
	.w2(32'h3ccc7130),
	.w3(32'hbba5c9c2),
	.w4(32'hbb80c565),
	.w5(32'hbb778019),
	.w6(32'h3c96d684),
	.w7(32'h3bef090c),
	.w8(32'hbbf3b921),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba26cf2d),
	.w1(32'h395976fd),
	.w2(32'h3d706443),
	.w3(32'h3c20a2b3),
	.w4(32'h3b0e00ad),
	.w5(32'hbbd762bf),
	.w6(32'hbc2ae007),
	.w7(32'hbc00f56c),
	.w8(32'hbb4628f2),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a141e37),
	.w1(32'h3ade9ed6),
	.w2(32'hbbd7bfdc),
	.w3(32'hbc7788d5),
	.w4(32'hbc0bf5b0),
	.w5(32'h3b42c29e),
	.w6(32'h3bf6b72c),
	.w7(32'h3d0e1df8),
	.w8(32'h3bb8f508),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae75fac),
	.w1(32'hbba46c58),
	.w2(32'h3b48d955),
	.w3(32'hbb3689e0),
	.w4(32'h3a81444d),
	.w5(32'h3b965bb8),
	.w6(32'hb97d06cc),
	.w7(32'hbb18751e),
	.w8(32'h3c8f7ebe),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe57bfd),
	.w1(32'hba58af1b),
	.w2(32'hbb6169a2),
	.w3(32'hbba10a42),
	.w4(32'hbb0007d2),
	.w5(32'hbb810b0a),
	.w6(32'h3ad72be6),
	.w7(32'h3ca18bb8),
	.w8(32'h3a760264),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf29dc6),
	.w1(32'h3a5df510),
	.w2(32'h3b2dbf33),
	.w3(32'h3b84d401),
	.w4(32'hbbb6e576),
	.w5(32'hbb24f6c0),
	.w6(32'hbbc386a5),
	.w7(32'hbb49ad8d),
	.w8(32'h3aecb1ce),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b48e087),
	.w1(32'hbbd3ef53),
	.w2(32'hba953aa3),
	.w3(32'hbc2fab6d),
	.w4(32'h3bdcbe0f),
	.w5(32'h3abb4a4c),
	.w6(32'h3a8f4a06),
	.w7(32'hba8285ca),
	.w8(32'h3968456c),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39283760),
	.w1(32'hbb06e090),
	.w2(32'h39997043),
	.w3(32'h3c5beee3),
	.w4(32'h397b2eb1),
	.w5(32'hba6f14b2),
	.w6(32'hba9a0d44),
	.w7(32'hbc3230e1),
	.w8(32'hbc054a9d),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1703c2),
	.w1(32'h3b0c047a),
	.w2(32'h3a6fec77),
	.w3(32'h3c3d9565),
	.w4(32'hbaf905a3),
	.w5(32'hba8c0562),
	.w6(32'hbb17a403),
	.w7(32'h3b38cf2f),
	.w8(32'h3ad3d59a),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba39798),
	.w1(32'h3aafb6ac),
	.w2(32'hb99388d2),
	.w3(32'hbb360318),
	.w4(32'h3b73487c),
	.w5(32'h3c2ed401),
	.w6(32'h3b6e4f21),
	.w7(32'hbaba533e),
	.w8(32'hbc396db0),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2f7038),
	.w1(32'hbbaa2949),
	.w2(32'h39509884),
	.w3(32'hbbb1a2cc),
	.w4(32'hbbdf29b1),
	.w5(32'h3c0b1967),
	.w6(32'h3a9b9ae3),
	.w7(32'h38fcce0f),
	.w8(32'h3b48411e),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaae552b),
	.w1(32'hbbc92313),
	.w2(32'h3c7d4440),
	.w3(32'h3bf6603b),
	.w4(32'h3b026adb),
	.w5(32'hba7879e8),
	.w6(32'h3ad2a7b7),
	.w7(32'h3c08e791),
	.w8(32'hbadd59de),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b86fdf8),
	.w1(32'hbb89dac5),
	.w2(32'hbbc5e4f9),
	.w3(32'hbb1930d5),
	.w4(32'hbb500f08),
	.w5(32'h3a385e65),
	.w6(32'h3b8db127),
	.w7(32'h38de7b15),
	.w8(32'hbbaec245),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9816ecc),
	.w1(32'hbab4af76),
	.w2(32'hbaa12582),
	.w3(32'h3afc524e),
	.w4(32'hbb0563c8),
	.w5(32'hba9005d3),
	.w6(32'h3a863a9d),
	.w7(32'h3a5b31c0),
	.w8(32'h39fd271e),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394fe431),
	.w1(32'h389f2cdf),
	.w2(32'h3ac10aa2),
	.w3(32'hbbbd2165),
	.w4(32'h384d1e6f),
	.w5(32'h3c6d6776),
	.w6(32'hbb98c001),
	.w7(32'hbb993f87),
	.w8(32'h3c466bf9),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9cd50a),
	.w1(32'h3ad042fc),
	.w2(32'h3adc71d5),
	.w3(32'hbc5cc3e4),
	.w4(32'hbc08ed40),
	.w5(32'hbc34e555),
	.w6(32'hba27dfb3),
	.w7(32'hba7efe35),
	.w8(32'hbbb5e5ca),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5d3939),
	.w1(32'hb9cab611),
	.w2(32'h3b597e30),
	.w3(32'h3b9f5dcb),
	.w4(32'h3bd81c41),
	.w5(32'h3b242182),
	.w6(32'h3a858ffc),
	.w7(32'h3aa8b89a),
	.w8(32'hba1c68cc),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb77956e),
	.w1(32'h3ba9d25d),
	.w2(32'h3c75cf0b),
	.w3(32'h3d623570),
	.w4(32'h3c0893c2),
	.w5(32'h3c613153),
	.w6(32'h3a457e72),
	.w7(32'hbc827380),
	.w8(32'h3c37b107),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afec9d6),
	.w1(32'hbcb8ea6e),
	.w2(32'h3b4652e3),
	.w3(32'h3da2cd42),
	.w4(32'h3b9f6c24),
	.w5(32'h3d330038),
	.w6(32'hbb9993d7),
	.w7(32'h3b508534),
	.w8(32'h3a85d17a),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae1f268),
	.w1(32'h3cf5475e),
	.w2(32'h3c04829e),
	.w3(32'h3c1199f4),
	.w4(32'hba9452ce),
	.w5(32'h39d082fe),
	.w6(32'h3bc85fa4),
	.w7(32'hb99df372),
	.w8(32'hbc33f951),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae5215f),
	.w1(32'hbd9173a5),
	.w2(32'hbcd14140),
	.w3(32'h39b429a8),
	.w4(32'h3c0329c1),
	.w5(32'hbc1180fc),
	.w6(32'hbbd7cb1d),
	.w7(32'hbd2214c3),
	.w8(32'h3b733519),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb17952),
	.w1(32'h3d074846),
	.w2(32'hbc0f9714),
	.w3(32'h3b18d7ab),
	.w4(32'h3b5720b5),
	.w5(32'hbd7c0ebb),
	.w6(32'h3b4771bb),
	.w7(32'h3bad9cf4),
	.w8(32'hbc74502c),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baa15ae),
	.w1(32'hbc834cf9),
	.w2(32'h390f8989),
	.w3(32'hba8ac0b2),
	.w4(32'hba08da7a),
	.w5(32'hbc50f62f),
	.w6(32'h392fb025),
	.w7(32'hbafed403),
	.w8(32'h3a191f8d),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c336759),
	.w1(32'hbb910e5c),
	.w2(32'hbc2176aa),
	.w3(32'h3afcac00),
	.w4(32'h3afffc34),
	.w5(32'hba746494),
	.w6(32'hbbc7d206),
	.w7(32'h3b2712fe),
	.w8(32'h3afd5f76),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d6946f2),
	.w1(32'hbd087978),
	.w2(32'hbc40e379),
	.w3(32'hbcdae9bc),
	.w4(32'h3b125674),
	.w5(32'h3b0c9a4f),
	.w6(32'hbc4d2310),
	.w7(32'hba18fb51),
	.w8(32'hbc453b0c),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d82f182),
	.w1(32'h3c911523),
	.w2(32'h3b7557f6),
	.w3(32'hbb4e3bbf),
	.w4(32'h3be5eeb0),
	.w5(32'h3b7fa0a3),
	.w6(32'hba2afe3d),
	.w7(32'hbc40e9ad),
	.w8(32'h3c03cfe3),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb38bac1),
	.w1(32'h39922b47),
	.w2(32'h3b22644c),
	.w3(32'hbc0ab90d),
	.w4(32'hbbbe3b58),
	.w5(32'h3b61c8a1),
	.w6(32'hbb70fdd2),
	.w7(32'hbbe44664),
	.w8(32'hbd8cea09),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8a4737),
	.w1(32'h3b2b8774),
	.w2(32'hbb82b997),
	.w3(32'h3b80fcca),
	.w4(32'hbc81bd00),
	.w5(32'h3b535555),
	.w6(32'hbb56a438),
	.w7(32'hbc97a15e),
	.w8(32'h3c216910),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9cab24),
	.w1(32'h3b38c515),
	.w2(32'hbb3752aa),
	.w3(32'h3b4ed8ee),
	.w4(32'h3c0613f4),
	.w5(32'h3a8e1fc7),
	.w6(32'h3c05affa),
	.w7(32'hb8a1da81),
	.w8(32'hbc24297b),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c31fecd),
	.w1(32'hbc82bf83),
	.w2(32'h3bbe076f),
	.w3(32'h3c2f8123),
	.w4(32'hba3194bc),
	.w5(32'h3bde907a),
	.w6(32'hbbf2d987),
	.w7(32'hbca965a3),
	.w8(32'hbc348931),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4d9671),
	.w1(32'h3b24b175),
	.w2(32'h3afd806a),
	.w3(32'h3c4fb9aa),
	.w4(32'h3b4a67fa),
	.w5(32'hbc42ad56),
	.w6(32'h3b95349e),
	.w7(32'hb9fe297a),
	.w8(32'h3b55fd0b),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc04645c),
	.w1(32'h3a53113d),
	.w2(32'hb9f9075d),
	.w3(32'hbb3c8000),
	.w4(32'hbaacef52),
	.w5(32'h39a32cd4),
	.w6(32'hbaece6fc),
	.w7(32'h3beb381c),
	.w8(32'h3b936f21),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbb59b9),
	.w1(32'h3c62e7e5),
	.w2(32'hba83cf28),
	.w3(32'h3ad1cc8f),
	.w4(32'hbb5abaf8),
	.w5(32'h3c1b9300),
	.w6(32'hbb24594e),
	.w7(32'h3b9302b2),
	.w8(32'hba408c24),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule