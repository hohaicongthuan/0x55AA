module layer_10_featuremap_400(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafde4c1),
	.w1(32'h3bc4bfd4),
	.w2(32'hb90288c0),
	.w3(32'hbbb07c80),
	.w4(32'h3bb937e6),
	.w5(32'hbc634717),
	.w6(32'h3aaba4a0),
	.w7(32'h3bc6a437),
	.w8(32'hba7c119a),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba65588c),
	.w1(32'hbab3d2e8),
	.w2(32'hbbd0e4fb),
	.w3(32'hbbdaee82),
	.w4(32'hbb8425ab),
	.w5(32'hbbc1f64b),
	.w6(32'hbafa4459),
	.w7(32'hbb5bc774),
	.w8(32'hbb7556c3),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad0f70b),
	.w1(32'h3b44d588),
	.w2(32'h3aa33d7a),
	.w3(32'h388b821f),
	.w4(32'hba9f731e),
	.w5(32'hbbe957a7),
	.w6(32'h3a989db5),
	.w7(32'hbbe3552d),
	.w8(32'hbac044dc),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7247d7),
	.w1(32'hbb1bd71f),
	.w2(32'hbadb92f2),
	.w3(32'h3bbdea92),
	.w4(32'hbc2a3663),
	.w5(32'hba4f5e36),
	.w6(32'h3b75f27f),
	.w7(32'hbc05bfdc),
	.w8(32'hbbcb8ebb),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2db1ee),
	.w1(32'hbbb443fa),
	.w2(32'h3b1cb6b5),
	.w3(32'hbbe3dd35),
	.w4(32'hbbcbc0ad),
	.w5(32'h3be0e4af),
	.w6(32'hba38ee8d),
	.w7(32'hbba39206),
	.w8(32'hb8a3ba1c),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6faab3),
	.w1(32'hbb1a7b15),
	.w2(32'hbac5fe5c),
	.w3(32'h3b93386a),
	.w4(32'hbb9fd4d8),
	.w5(32'h3a9862c7),
	.w6(32'hbaf44aff),
	.w7(32'h3b120ec8),
	.w8(32'hba9e5cfe),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbacef72a),
	.w1(32'hba9239ed),
	.w2(32'h3be89a46),
	.w3(32'hbb94525e),
	.w4(32'hbb2c88bd),
	.w5(32'h3c064d51),
	.w6(32'hbba61f07),
	.w7(32'h3b11fe87),
	.w8(32'h3bfb4fa0),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba003c0d),
	.w1(32'hbae9fc92),
	.w2(32'h3c23d6dd),
	.w3(32'hbbc5b603),
	.w4(32'h3b697e41),
	.w5(32'hbb8e3154),
	.w6(32'h3ba68225),
	.w7(32'h3bc209d5),
	.w8(32'h3b680c81),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaed7f2e),
	.w1(32'h3986b7c1),
	.w2(32'h3b1626a1),
	.w3(32'hbc11390b),
	.w4(32'hbb8c7aea),
	.w5(32'h3b289fc6),
	.w6(32'hbb92eb75),
	.w7(32'hbb5bb123),
	.w8(32'hba82d5a9),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbcb919),
	.w1(32'h3bc750f0),
	.w2(32'h3c2f8018),
	.w3(32'hbb738021),
	.w4(32'h3a93cc6a),
	.w5(32'h3b616a2e),
	.w6(32'hbbb35cee),
	.w7(32'hbbc8a9e2),
	.w8(32'hbbf64c98),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b82ed8b),
	.w1(32'h3abcfcac),
	.w2(32'h3bd1ca15),
	.w3(32'h3b08b4b0),
	.w4(32'h3b38787b),
	.w5(32'h3b50ec1e),
	.w6(32'hbb7d5ef1),
	.w7(32'h3a8ca353),
	.w8(32'h3acce1fa),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b69fa59),
	.w1(32'hbbd676de),
	.w2(32'h3c0adaaf),
	.w3(32'h3b799232),
	.w4(32'hbbbc6c75),
	.w5(32'h3c990083),
	.w6(32'h3a727b6b),
	.w7(32'hb9e289f9),
	.w8(32'h3c20e0e4),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4ed3cf),
	.w1(32'h3b174834),
	.w2(32'h3b7f0a4a),
	.w3(32'h3bffcc94),
	.w4(32'hbc218cbf),
	.w5(32'h3c5ea45f),
	.w6(32'hbb8a52a0),
	.w7(32'hbc2e814c),
	.w8(32'hbb45cd7b),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd9fa0b),
	.w1(32'hbac9e924),
	.w2(32'h3b0e8105),
	.w3(32'hbb8e0ce0),
	.w4(32'h3b33c437),
	.w5(32'hbba5eb64),
	.w6(32'hbbab3ce8),
	.w7(32'hb7b6148e),
	.w8(32'h39a408d7),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38a60858),
	.w1(32'hbbabb713),
	.w2(32'hbc46db85),
	.w3(32'hbaef11c5),
	.w4(32'hbb8909ac),
	.w5(32'hbb3ad764),
	.w6(32'hbb8ebf93),
	.w7(32'hbb61f0bc),
	.w8(32'hbc08f5aa),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb774ff4),
	.w1(32'hbb75182d),
	.w2(32'hbbfd26f9),
	.w3(32'hbbbd5d58),
	.w4(32'hbac74705),
	.w5(32'h3bd94c73),
	.w6(32'hbc112d93),
	.w7(32'hbadddcce),
	.w8(32'h3a605cef),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2c69bb),
	.w1(32'hb99e55d5),
	.w2(32'hbaae8eed),
	.w3(32'hbbfec1dc),
	.w4(32'hbb4fc1c9),
	.w5(32'h3b286133),
	.w6(32'hbbd97d1c),
	.w7(32'hbb864f2b),
	.w8(32'hba381740),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a386940),
	.w1(32'h3cac341f),
	.w2(32'h3cf63953),
	.w3(32'h3b4a3d66),
	.w4(32'h3c412b25),
	.w5(32'h3bd6d71f),
	.w6(32'h3b9857a8),
	.w7(32'h3c8b5cf2),
	.w8(32'h3c119eef),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a56e3cd),
	.w1(32'hbb925548),
	.w2(32'h3b99dff2),
	.w3(32'hbbdf8e08),
	.w4(32'hbc0d3a5e),
	.w5(32'h3c8a8f80),
	.w6(32'h3b14237f),
	.w7(32'hbbbaa0eb),
	.w8(32'h3b01d517),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba02d8d),
	.w1(32'hbc15d424),
	.w2(32'hbbe5ac91),
	.w3(32'hbb309c9b),
	.w4(32'hbbbf1fe5),
	.w5(32'hbbd65c2d),
	.w6(32'hbc0f2460),
	.w7(32'hbb02b38a),
	.w8(32'hbbfaba16),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc25be9a),
	.w1(32'hb9a03749),
	.w2(32'h3bfc0db5),
	.w3(32'hbc4bb800),
	.w4(32'h39a59dee),
	.w5(32'h3c84161c),
	.w6(32'hbc200dae),
	.w7(32'h3b60e631),
	.w8(32'h3c0c3f15),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9f71f2),
	.w1(32'h3b0678f7),
	.w2(32'hba6841b4),
	.w3(32'h3c12b95b),
	.w4(32'hbaa5b288),
	.w5(32'h3b362e5f),
	.w6(32'h3b2e63af),
	.w7(32'h3b8f6377),
	.w8(32'h3ae7d6db),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b78286b),
	.w1(32'h3c0e8a5a),
	.w2(32'h3c553f10),
	.w3(32'hbbc1a215),
	.w4(32'hbb54e84c),
	.w5(32'h3c4417f2),
	.w6(32'h3b9df105),
	.w7(32'h3c6851a7),
	.w8(32'h3b78028b),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1b1119),
	.w1(32'h3a0c5c01),
	.w2(32'hbb4cbbb5),
	.w3(32'h3bac0968),
	.w4(32'h3b82f0fd),
	.w5(32'h3ab80748),
	.w6(32'hbb55c3ed),
	.w7(32'hbbd1e068),
	.w8(32'hbbf1b710),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf5adda),
	.w1(32'hbb24aed7),
	.w2(32'hbb5b683e),
	.w3(32'h3bf4253d),
	.w4(32'hbb3dd324),
	.w5(32'hbbe56d6f),
	.w6(32'h3ad20118),
	.w7(32'h3a17c93c),
	.w8(32'hbb5d89f0),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad86281),
	.w1(32'h3879cf27),
	.w2(32'h3ba51e90),
	.w3(32'hbbcb2533),
	.w4(32'hbaee6603),
	.w5(32'h3b831c3a),
	.w6(32'hbc03781a),
	.w7(32'h3b002e5f),
	.w8(32'h3b8b3e76),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b39cf0d),
	.w1(32'hbada6736),
	.w2(32'hbb2a22bc),
	.w3(32'h38bd391b),
	.w4(32'hbba21d9f),
	.w5(32'hbb3a9065),
	.w6(32'h3b1b402f),
	.w7(32'hbaadbf9b),
	.w8(32'h3b7166c6),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac094bb),
	.w1(32'h3b6c9328),
	.w2(32'h3b912775),
	.w3(32'hbadcb47d),
	.w4(32'h3b877b05),
	.w5(32'h3a978bcc),
	.w6(32'hbb504c6b),
	.w7(32'h3b2839be),
	.w8(32'hbb20e5a9),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a784076),
	.w1(32'hbbb87e4d),
	.w2(32'hba7e2643),
	.w3(32'hbb0a26cb),
	.w4(32'hb9f9cdf1),
	.w5(32'h393dcc67),
	.w6(32'h3a878883),
	.w7(32'hbaf5ec66),
	.w8(32'hb9867ec7),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4c524c),
	.w1(32'hbb228dc8),
	.w2(32'h3b870d3a),
	.w3(32'h3adb388f),
	.w4(32'hbb8af149),
	.w5(32'h3c09fc2f),
	.w6(32'hbb9a89c2),
	.w7(32'h392d5bb8),
	.w8(32'h3a9ec3ce),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1b0928),
	.w1(32'hbaeb0212),
	.w2(32'hbaeee1c6),
	.w3(32'h3c5d60da),
	.w4(32'hbbadd3cc),
	.w5(32'hbb4e26bd),
	.w6(32'h3bf43317),
	.w7(32'hbad93107),
	.w8(32'h3afe4624),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3192b2),
	.w1(32'hba22b9cb),
	.w2(32'hbb34d00e),
	.w3(32'h3bd7392b),
	.w4(32'h3aeb0bbb),
	.w5(32'hbb0abee4),
	.w6(32'h3be925ea),
	.w7(32'hbbb6c177),
	.w8(32'hbbbb06d8),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a69d4ac),
	.w1(32'hba517810),
	.w2(32'h3a662b57),
	.w3(32'h3b203acd),
	.w4(32'hbaedd030),
	.w5(32'h390e69c1),
	.w6(32'h3af865ce),
	.w7(32'hbb25e28b),
	.w8(32'hba71e7ac),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ccb8a1),
	.w1(32'h3b2d1407),
	.w2(32'h3aa25e4d),
	.w3(32'hba39fcba),
	.w4(32'hbb3fb61f),
	.w5(32'hbbadac15),
	.w6(32'hbb2d4594),
	.w7(32'hbbaac0ab),
	.w8(32'hbc14d963),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba33fe9b),
	.w1(32'h3a83ea2e),
	.w2(32'h3c13c736),
	.w3(32'hbbc8d446),
	.w4(32'hba56763c),
	.w5(32'h3a19fdda),
	.w6(32'hbc01b3e8),
	.w7(32'h3b539257),
	.w8(32'h3bf3f6b4),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bea52bc),
	.w1(32'h3bb50ee8),
	.w2(32'h3c062a81),
	.w3(32'hbaa75a8a),
	.w4(32'h3be638b2),
	.w5(32'h3b370904),
	.w6(32'h3bf91f51),
	.w7(32'hb780e96a),
	.w8(32'h3b3c9548),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adbeed6),
	.w1(32'hbc82ac2c),
	.w2(32'hbbac42a1),
	.w3(32'hbbaa571f),
	.w4(32'hbc51a540),
	.w5(32'hbb46ea32),
	.w6(32'h3b190c16),
	.w7(32'hbc158cfd),
	.w8(32'hbb887baf),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfbc348),
	.w1(32'h3b55926b),
	.w2(32'hbc5ec9fd),
	.w3(32'h39b1d3a8),
	.w4(32'h3a9c809e),
	.w5(32'hbb3497c5),
	.w6(32'h39326e16),
	.w7(32'h3b944742),
	.w8(32'h3b393874),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc328ee),
	.w1(32'h3c385b06),
	.w2(32'hbc14a4e0),
	.w3(32'h3b807568),
	.w4(32'h3c3f4653),
	.w5(32'hbc7b14a5),
	.w6(32'h3b74eb0d),
	.w7(32'h3c43410a),
	.w8(32'hbb8372db),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6bb90e),
	.w1(32'hbbbb8093),
	.w2(32'hbc0c85d4),
	.w3(32'hbc0a8495),
	.w4(32'hbb580c4e),
	.w5(32'hbbf8ec59),
	.w6(32'hbb9bb102),
	.w7(32'hbc00d2be),
	.w8(32'hbbfff437),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaef823d),
	.w1(32'hb9fc11bd),
	.w2(32'hb98ce67f),
	.w3(32'hbaab73f8),
	.w4(32'hb8c5da33),
	.w5(32'h3b18d4be),
	.w6(32'hbb693258),
	.w7(32'h3aad62d7),
	.w8(32'hba751b72),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3997f347),
	.w1(32'hbb33a729),
	.w2(32'hbb5bd624),
	.w3(32'h3bd3245d),
	.w4(32'hbb873f74),
	.w5(32'h3bdb01a7),
	.w6(32'h3b00f4cf),
	.w7(32'hbaa3c3f5),
	.w8(32'hbba98432),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8bee31),
	.w1(32'hbaf2d582),
	.w2(32'hbb640ae1),
	.w3(32'h3bb6d0c6),
	.w4(32'hbbf5e2b2),
	.w5(32'h3ba6b986),
	.w6(32'hb973d258),
	.w7(32'hbbb9946b),
	.w8(32'hbb90653e),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b008069),
	.w1(32'h3bf66985),
	.w2(32'h3be0e163),
	.w3(32'hbaebb8c4),
	.w4(32'h3c278ff0),
	.w5(32'hbc6a2bf4),
	.w6(32'hbb94519a),
	.w7(32'h3bc4bd57),
	.w8(32'hbc154473),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bace63c),
	.w1(32'h3af4821d),
	.w2(32'hbb6357b5),
	.w3(32'h3b2e8ca3),
	.w4(32'hb78df0d6),
	.w5(32'hb98b80a0),
	.w6(32'h38f3d80d),
	.w7(32'hba9945ac),
	.w8(32'hbc0a8299),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a71377),
	.w1(32'h3a858773),
	.w2(32'hbbd7f698),
	.w3(32'hbb64a776),
	.w4(32'hb8b9e549),
	.w5(32'hbbbbfc64),
	.w6(32'hbb8d17ba),
	.w7(32'hbbb460c0),
	.w8(32'hbb5e31a5),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9ff73d),
	.w1(32'hbad6306b),
	.w2(32'hbc075ff4),
	.w3(32'h3ab1d1b4),
	.w4(32'hbb61d9aa),
	.w5(32'hbc471009),
	.w6(32'h3b3e3d76),
	.w7(32'h398a1dbe),
	.w8(32'hbb845b70),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf42713),
	.w1(32'h3c08d5b1),
	.w2(32'h3c9eb76f),
	.w3(32'hbc680d8c),
	.w4(32'hba7887b1),
	.w5(32'h3c1e9ffa),
	.w6(32'hbba16451),
	.w7(32'hba809218),
	.w8(32'h3b4e4562),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb18780c),
	.w1(32'h3ace8426),
	.w2(32'h3b9261e1),
	.w3(32'hbbd22735),
	.w4(32'h3c11502a),
	.w5(32'h3b050869),
	.w6(32'hbb82ec61),
	.w7(32'h3c1dcfc0),
	.w8(32'h3bfa9958),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3a9194),
	.w1(32'h3b1b5859),
	.w2(32'h3bb2bfc5),
	.w3(32'hbb66de5a),
	.w4(32'h3c68225f),
	.w5(32'h3b0c1ad8),
	.w6(32'hbbd1e9ca),
	.w7(32'h3b286ef8),
	.w8(32'h3a8caeab),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b11abd8),
	.w1(32'h3a73d8cc),
	.w2(32'hbb1926fe),
	.w3(32'h3bd17332),
	.w4(32'h3b44633a),
	.w5(32'h3b883763),
	.w6(32'h3ab0768a),
	.w7(32'hbb9955ea),
	.w8(32'h3a6b1650),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b624fa9),
	.w1(32'hbaf2ea0a),
	.w2(32'hb8e59820),
	.w3(32'h3ca7a51c),
	.w4(32'hbc368c5b),
	.w5(32'hbab38ff7),
	.w6(32'h3b5280c9),
	.w7(32'hbb94e0d0),
	.w8(32'hbaf513a2),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9bafb55),
	.w1(32'h3b57515c),
	.w2(32'h3bd88622),
	.w3(32'hbb3382a2),
	.w4(32'h3b488445),
	.w5(32'hbb183361),
	.w6(32'hbb225c65),
	.w7(32'h3b59aac9),
	.w8(32'h399ed4b6),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf11b77),
	.w1(32'h3c10c8ca),
	.w2(32'h3cb2cbd5),
	.w3(32'hbb2b39df),
	.w4(32'h3b150799),
	.w5(32'h3c36a3c9),
	.w6(32'h39ed665d),
	.w7(32'hbaa83212),
	.w8(32'h3b9398bf),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b97ec2c),
	.w1(32'h3b34eb5a),
	.w2(32'h3af3613d),
	.w3(32'hbac362a1),
	.w4(32'h3b85b25f),
	.w5(32'h3bbb078f),
	.w6(32'hba42a550),
	.w7(32'hba8f86a3),
	.w8(32'h3b1432d9),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3b2103),
	.w1(32'hbb85320c),
	.w2(32'hbbca57fe),
	.w3(32'hba99fd8b),
	.w4(32'hbbf054d6),
	.w5(32'hbbc1d651),
	.w6(32'h39ae6d44),
	.w7(32'hbbdf0ecd),
	.w8(32'hbb34759f),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0b23eb),
	.w1(32'hbbf87bf3),
	.w2(32'hbab5201f),
	.w3(32'hbb0298ce),
	.w4(32'hbc93325c),
	.w5(32'h3c8900f4),
	.w6(32'hbb941747),
	.w7(32'hbc37f54b),
	.w8(32'h3b2fcfad),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a32d86f),
	.w1(32'hbb314423),
	.w2(32'hbb60d452),
	.w3(32'h3bb388e7),
	.w4(32'hbacd5cd7),
	.w5(32'hbae0c00d),
	.w6(32'hb829b270),
	.w7(32'hb99a4026),
	.w8(32'hbbe43656),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f48d8),
	.w1(32'h3c1b4046),
	.w2(32'hbbdd4311),
	.w3(32'hbb93997b),
	.w4(32'h3b7eb452),
	.w5(32'hbb26c4f6),
	.w6(32'hbc129461),
	.w7(32'h3b5c280b),
	.w8(32'hba8fe838),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba56bbf),
	.w1(32'hbc4885a8),
	.w2(32'hbbdb960e),
	.w3(32'h3b8b76a2),
	.w4(32'hbb056766),
	.w5(32'hbb8c6822),
	.w6(32'h3b74fda6),
	.w7(32'hbbc1cd66),
	.w8(32'h3b3c7477),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba95502),
	.w1(32'h3a406a34),
	.w2(32'h3c1de26e),
	.w3(32'hb8785610),
	.w4(32'h3a0b7395),
	.w5(32'h3c0e6af6),
	.w6(32'hbba8b2d5),
	.w7(32'hba69a695),
	.w8(32'h3b86a5e7),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a93962c),
	.w1(32'h3ab46014),
	.w2(32'h3bd4890c),
	.w3(32'hb9aa1d3d),
	.w4(32'h3ac5ffd2),
	.w5(32'h3c48707b),
	.w6(32'h3ac50d51),
	.w7(32'h3b43530c),
	.w8(32'h3c219d74),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b22042c),
	.w1(32'hbb27aef6),
	.w2(32'hbbe7ae6f),
	.w3(32'h3a74e6fa),
	.w4(32'h3b4da4c2),
	.w5(32'hbbf7adf0),
	.w6(32'h3a3a7dc0),
	.w7(32'hbb8cb60e),
	.w8(32'hbc065d9e),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe6a3ef),
	.w1(32'hbc475aac),
	.w2(32'hbae7d4cd),
	.w3(32'hbbc0f86f),
	.w4(32'hbc7a024d),
	.w5(32'h3c35474e),
	.w6(32'hbb136757),
	.w7(32'hbb7f6ec7),
	.w8(32'h3bc5f5c0),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad6a1b9),
	.w1(32'h3b194e2b),
	.w2(32'h3bb07b52),
	.w3(32'h3be11df2),
	.w4(32'h3a957f0f),
	.w5(32'h3b84f068),
	.w6(32'hba1cd531),
	.w7(32'hbaf2a5e3),
	.w8(32'h3b1653aa),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1f4046),
	.w1(32'hba6f2d96),
	.w2(32'h3ae08501),
	.w3(32'h38ece951),
	.w4(32'hb9dff354),
	.w5(32'h3b538264),
	.w6(32'hbb627a5f),
	.w7(32'h3b7027c3),
	.w8(32'h3b63f4bd),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e6a34),
	.w1(32'h3a3a2a2f),
	.w2(32'h3c022d85),
	.w3(32'hbc225c6b),
	.w4(32'hbb1b21c6),
	.w5(32'h3bc67289),
	.w6(32'hbbded79d),
	.w7(32'hbc2a8dc9),
	.w8(32'h3a22d97a),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb0c7dd),
	.w1(32'h3be2fc38),
	.w2(32'h3c3a6743),
	.w3(32'h3a96cc7d),
	.w4(32'h3c47f7a5),
	.w5(32'h3c35eb5e),
	.w6(32'h3abad267),
	.w7(32'h3b04a4fd),
	.w8(32'h3bd76c99),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a071164),
	.w1(32'h3b389c6c),
	.w2(32'h3c0308c2),
	.w3(32'hbaee176b),
	.w4(32'h3c2aa3d6),
	.w5(32'h3bfdd09e),
	.w6(32'h3bee9409),
	.w7(32'h3c4bdec0),
	.w8(32'h3c89c485),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1271e9),
	.w1(32'h3af5d4d3),
	.w2(32'h3a15b71e),
	.w3(32'h3bcaf3eb),
	.w4(32'hbb631fb4),
	.w5(32'hbc425b8a),
	.w6(32'h3c46d15f),
	.w7(32'h3c3222a1),
	.w8(32'hbc35c060),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b932232),
	.w1(32'hbbfb051d),
	.w2(32'h3abfa2ed),
	.w3(32'h3a1d90e9),
	.w4(32'hba3d1ba4),
	.w5(32'hbb2e4605),
	.w6(32'hbbe981aa),
	.w7(32'hbb970ddb),
	.w8(32'hbacafb32),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bacd2dd),
	.w1(32'hbaa3ef91),
	.w2(32'h3b28c3b8),
	.w3(32'h3a590b81),
	.w4(32'h39f559b1),
	.w5(32'h3a0a61a7),
	.w6(32'hbb19133f),
	.w7(32'h3ba0402c),
	.w8(32'h3c31ff7b),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbad623a),
	.w1(32'hbb82ef1a),
	.w2(32'hbbd0f63a),
	.w3(32'hbbff54cb),
	.w4(32'h3b19a66e),
	.w5(32'h3ac2bad6),
	.w6(32'h3aebafae),
	.w7(32'h3c741522),
	.w8(32'h3bbea7c6),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4ac36f),
	.w1(32'hbb8af790),
	.w2(32'h3b8d118c),
	.w3(32'hb9e868d9),
	.w4(32'h3bb30530),
	.w5(32'h3b7fa2d4),
	.w6(32'h3b3dcdf8),
	.w7(32'h3b954e57),
	.w8(32'h3bc58929),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b108d25),
	.w1(32'h3b1031a6),
	.w2(32'h3c22c805),
	.w3(32'h3a9fbbbc),
	.w4(32'h3bd1d811),
	.w5(32'h3d0c8a16),
	.w6(32'hbba55e09),
	.w7(32'hbc33f66b),
	.w8(32'hbba73ffa),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2884fb),
	.w1(32'h3916fb9e),
	.w2(32'h3b61c6ce),
	.w3(32'h3bd5645e),
	.w4(32'h3ae95b43),
	.w5(32'h3c0a348b),
	.w6(32'hbb569e6f),
	.w7(32'h3b4f13e5),
	.w8(32'h3bfc3cdc),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc4335ec),
	.w1(32'hbbfbd4f8),
	.w2(32'h3b29c19a),
	.w3(32'hbbafbfc9),
	.w4(32'h3b45727b),
	.w5(32'hbaa461bb),
	.w6(32'h3b1011a1),
	.w7(32'h3b88e0f4),
	.w8(32'h3c952014),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6d958f),
	.w1(32'hba549447),
	.w2(32'h3b76c76b),
	.w3(32'hbbc7dd32),
	.w4(32'hbc2f57e8),
	.w5(32'hbb6f779d),
	.w6(32'hbbc0b56b),
	.w7(32'hbc25c1cf),
	.w8(32'hbbdbd46a),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c240542),
	.w1(32'hbb16c7e4),
	.w2(32'h3ada453e),
	.w3(32'h3a9d4775),
	.w4(32'h3b8d29a8),
	.w5(32'h3b6e2210),
	.w6(32'hbadf36db),
	.w7(32'h3c2a117e),
	.w8(32'h3c2ff409),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba9c3d1),
	.w1(32'hb655d334),
	.w2(32'h3c6e9054),
	.w3(32'hba33172d),
	.w4(32'h3c2eb896),
	.w5(32'h3c99c9d0),
	.w6(32'hbb1feb0a),
	.w7(32'hbabeed83),
	.w8(32'h3aab09ad),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba56bfa),
	.w1(32'h3bda18c0),
	.w2(32'h37e47630),
	.w3(32'h3bcf77f8),
	.w4(32'h3c31c744),
	.w5(32'h3a032b1c),
	.w6(32'h3b224126),
	.w7(32'h3c91f010),
	.w8(32'h3c65983c),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2209a4),
	.w1(32'hbb433e4c),
	.w2(32'h3b2c800e),
	.w3(32'h3c108f03),
	.w4(32'h3ab42d1f),
	.w5(32'h39418c62),
	.w6(32'h3b936366),
	.w7(32'h3b8af7dc),
	.w8(32'h3ba20abf),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba91127f),
	.w1(32'hbb7487db),
	.w2(32'hbb597dc0),
	.w3(32'hbb22431c),
	.w4(32'h3b1e857e),
	.w5(32'hba78f5a3),
	.w6(32'hb9e00142),
	.w7(32'hbae1fb57),
	.w8(32'hba8e6265),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb452977),
	.w1(32'hb99872b3),
	.w2(32'h3a0bab4a),
	.w3(32'h39634053),
	.w4(32'h3c485e66),
	.w5(32'h3bb98b74),
	.w6(32'hbb9d2bf9),
	.w7(32'h3c1bda0d),
	.w8(32'h3b95220c),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2564e6),
	.w1(32'hbbe54203),
	.w2(32'hbbe3a333),
	.w3(32'h3ba26061),
	.w4(32'hbb07f521),
	.w5(32'hbb398986),
	.w6(32'hba5fcd19),
	.w7(32'h3bd51099),
	.w8(32'h3bbe8857),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb92e6b4),
	.w1(32'h3a67ea48),
	.w2(32'hba70885b),
	.w3(32'hbb3bebc7),
	.w4(32'hba9517c3),
	.w5(32'hbc22ff6b),
	.w6(32'h3b975bbf),
	.w7(32'hbbab8e6a),
	.w8(32'hbbce52aa),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1fb94d),
	.w1(32'hbb703eac),
	.w2(32'hbbe6168a),
	.w3(32'hbc27913d),
	.w4(32'h3a85066d),
	.w5(32'h3ab42800),
	.w6(32'hbba40351),
	.w7(32'h3a7f3410),
	.w8(32'hbb964b47),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3457f6),
	.w1(32'hba2becbb),
	.w2(32'hbb425e53),
	.w3(32'hbb8b65b8),
	.w4(32'hbadfadff),
	.w5(32'hb9e98e98),
	.w6(32'hbb91ab32),
	.w7(32'h39f5c760),
	.w8(32'h3b7b47f2),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaec4eaa),
	.w1(32'hba08f8a5),
	.w2(32'hbb1f9a0d),
	.w3(32'hbb7af94f),
	.w4(32'hba2a812e),
	.w5(32'hbba8a107),
	.w6(32'h3aa043e8),
	.w7(32'hba0bfb78),
	.w8(32'h3b4c8cf2),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af55a5c),
	.w1(32'h3bd1e88f),
	.w2(32'h3bc4e115),
	.w3(32'hba9a8dfc),
	.w4(32'h3bdd8ca4),
	.w5(32'h3c296de6),
	.w6(32'h3b5d9ac3),
	.w7(32'hb99667b6),
	.w8(32'h3ca51a30),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1331f2),
	.w1(32'hbc2ccf83),
	.w2(32'hbc709fe3),
	.w3(32'h3a97f3b7),
	.w4(32'hbb413410),
	.w5(32'hbbec82f2),
	.w6(32'h3baef431),
	.w7(32'h394d9361),
	.w8(32'h3a63d867),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf3f364),
	.w1(32'hbaa7de67),
	.w2(32'h3c45420a),
	.w3(32'hbba52060),
	.w4(32'hbc247933),
	.w5(32'h3bb40641),
	.w6(32'hbc35295b),
	.w7(32'hbb862802),
	.w8(32'h3bcb5464),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b431c6a),
	.w1(32'hbc1bb870),
	.w2(32'hbc1e7dd5),
	.w3(32'h3b3aea18),
	.w4(32'hb7a3b550),
	.w5(32'hbc8753b4),
	.w6(32'hbacef70e),
	.w7(32'h3c84c34f),
	.w8(32'h3b87c4bc),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba416c0),
	.w1(32'hbb42697a),
	.w2(32'hbae9b1da),
	.w3(32'hbc25d87f),
	.w4(32'hbb393880),
	.w5(32'hbc621d29),
	.w6(32'hbac5f785),
	.w7(32'h3c104233),
	.w8(32'h3ba76774),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb141eb7),
	.w1(32'h39fcd4bf),
	.w2(32'h3a2929cd),
	.w3(32'hbba810f7),
	.w4(32'h3ca24a1c),
	.w5(32'h3cc25ecc),
	.w6(32'hbbff8e73),
	.w7(32'hb97d9972),
	.w8(32'h3bbf9654),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be3273f),
	.w1(32'h3b9efc53),
	.w2(32'h3ba5576d),
	.w3(32'hbac9a25e),
	.w4(32'hbb3946a9),
	.w5(32'hbc1ae599),
	.w6(32'h3b27bde3),
	.w7(32'hbb019e59),
	.w8(32'hbc22bb91),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad6a0a8),
	.w1(32'hbbacd4f2),
	.w2(32'hb9c38d7a),
	.w3(32'hbbd8e3f2),
	.w4(32'hba32340e),
	.w5(32'h3a05b734),
	.w6(32'hbb134d47),
	.w7(32'hbb26b1df),
	.w8(32'h3ab6e9b1),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1aa3f5),
	.w1(32'h3c423df7),
	.w2(32'h3c58ee8d),
	.w3(32'hbb54d4ee),
	.w4(32'h3c8fe445),
	.w5(32'h3c939897),
	.w6(32'h3b3fbc4a),
	.w7(32'h3b70377d),
	.w8(32'h3cc8952c),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae9f847),
	.w1(32'hbb0ab1ea),
	.w2(32'h3bc12d38),
	.w3(32'h3bc8499a),
	.w4(32'h3cd86756),
	.w5(32'h3cc64856),
	.w6(32'h3c15e090),
	.w7(32'h3cae1feb),
	.w8(32'h3d558c18),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92627fb),
	.w1(32'h3a2209dd),
	.w2(32'h3b9fdcd6),
	.w3(32'h3c9cc2d4),
	.w4(32'hbb0ab9b0),
	.w5(32'h3cb29141),
	.w6(32'h3ce74b0d),
	.w7(32'hbbb428ec),
	.w8(32'h38976808),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c487e28),
	.w1(32'hbb8011c2),
	.w2(32'hbc8b222b),
	.w3(32'h3b4fd092),
	.w4(32'h3c08d13d),
	.w5(32'h3a3b78d1),
	.w6(32'h3ac611c4),
	.w7(32'h3b9bc119),
	.w8(32'h3b808392),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb5ec11),
	.w1(32'h3a1ea83a),
	.w2(32'hbc0a3cad),
	.w3(32'h3bb57428),
	.w4(32'hbb07c6ab),
	.w5(32'hbb89051b),
	.w6(32'hbba70ff9),
	.w7(32'hba774a41),
	.w8(32'h39494f50),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb859968),
	.w1(32'h3ae3d0d9),
	.w2(32'h3c498999),
	.w3(32'hbb828245),
	.w4(32'h3bded5b8),
	.w5(32'h3c016d60),
	.w6(32'h3be30d8a),
	.w7(32'h3bccc37f),
	.w8(32'h3b9093e8),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9c42cf),
	.w1(32'h3b9b0728),
	.w2(32'h3b87a5cd),
	.w3(32'h3bd69e33),
	.w4(32'h3b6718b6),
	.w5(32'hba97a7b0),
	.w6(32'hbbb04ad1),
	.w7(32'h3c050fd1),
	.w8(32'h3bebcf6a),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf13a87),
	.w1(32'h3a850d66),
	.w2(32'h3c7df62d),
	.w3(32'h3ac96ae1),
	.w4(32'h3bf714d2),
	.w5(32'h3c192308),
	.w6(32'h3c6bf514),
	.w7(32'hbb7bc033),
	.w8(32'h3c34eaff),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc80ff4),
	.w1(32'h3b5b5b04),
	.w2(32'hbb5ba8e3),
	.w3(32'hbbf0fc12),
	.w4(32'h3be5b30c),
	.w5(32'hbb205e3b),
	.w6(32'hbac58296),
	.w7(32'hbab2859f),
	.w8(32'h3b884d1b),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa5b24d),
	.w1(32'hbb907de5),
	.w2(32'h3b07e2e7),
	.w3(32'hbb32f912),
	.w4(32'hbb4dad3d),
	.w5(32'hbb5dc4c8),
	.w6(32'hba10a755),
	.w7(32'hbc0cfdde),
	.w8(32'hbb6a6756),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8c3282),
	.w1(32'hbbc46879),
	.w2(32'hbb0ffadd),
	.w3(32'h3a287ae2),
	.w4(32'hbaf02300),
	.w5(32'h39e1b058),
	.w6(32'hbb5b103b),
	.w7(32'h3c376d9a),
	.w8(32'h3b61f0ec),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3e6e43),
	.w1(32'h3a3caccd),
	.w2(32'hbb620f3a),
	.w3(32'hbc0b8213),
	.w4(32'h3c0e2afe),
	.w5(32'h3bda843c),
	.w6(32'hbbfce637),
	.w7(32'hbbe7b58b),
	.w8(32'hbb0cbf60),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad7daf9),
	.w1(32'h3be3a649),
	.w2(32'h3c04fcd0),
	.w3(32'h3b0e25fd),
	.w4(32'hbaab4a03),
	.w5(32'h3ae38051),
	.w6(32'h3aeb0e28),
	.w7(32'hbbc3ba17),
	.w8(32'hbc221271),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b933684),
	.w1(32'h3b0a1924),
	.w2(32'hbb83e6b5),
	.w3(32'h38b5576e),
	.w4(32'hbb9443e9),
	.w5(32'hbbbbf0b0),
	.w6(32'h3ac67241),
	.w7(32'hb8b9bb14),
	.w8(32'hbae7d469),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf1f891),
	.w1(32'h3b69e819),
	.w2(32'hb9e577e7),
	.w3(32'hbb692c60),
	.w4(32'h3b6fe7e1),
	.w5(32'hba5024a5),
	.w6(32'h3b20e91f),
	.w7(32'hbb81bd25),
	.w8(32'h3c1c8253),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5c6d21),
	.w1(32'hbbcffd95),
	.w2(32'hbb9429c3),
	.w3(32'h38900f78),
	.w4(32'hbb94b8ee),
	.w5(32'h3b0301a5),
	.w6(32'h3b96735e),
	.w7(32'hbb122fee),
	.w8(32'h3a8c5c32),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6dc35e),
	.w1(32'hbba02f25),
	.w2(32'h3c118b3d),
	.w3(32'h3c4e87f1),
	.w4(32'hb8277519),
	.w5(32'h3ad75e7b),
	.w6(32'h38fed952),
	.w7(32'h3b5066d1),
	.w8(32'h3a9b2872),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b224c64),
	.w1(32'h3b1fe27f),
	.w2(32'h395530e3),
	.w3(32'hbb8ae2d2),
	.w4(32'hba83db5b),
	.w5(32'hbbcbeec3),
	.w6(32'hbba1b53f),
	.w7(32'h3bb1443d),
	.w8(32'hbb1e3970),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae19c81),
	.w1(32'hbb9a6321),
	.w2(32'hba081af1),
	.w3(32'hbb0a3f4c),
	.w4(32'h3b8e82b0),
	.w5(32'hbb4766eb),
	.w6(32'hba467327),
	.w7(32'h3c077ad1),
	.w8(32'h3b5c7707),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0dd1ba),
	.w1(32'h3b9090c1),
	.w2(32'hbbb70e90),
	.w3(32'h3a041dd2),
	.w4(32'h3b93c477),
	.w5(32'h3aaf5c69),
	.w6(32'h3afa3c27),
	.w7(32'h3b40e2a1),
	.w8(32'h39c65fa4),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b23f5fc),
	.w1(32'hbbb74021),
	.w2(32'h3b00795d),
	.w3(32'hbb47568e),
	.w4(32'h3b8f42cc),
	.w5(32'hbb107136),
	.w6(32'h3a964552),
	.w7(32'h3a776fc4),
	.w8(32'h3bc468d5),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1b8239),
	.w1(32'hbaaa766a),
	.w2(32'hbac82c17),
	.w3(32'h3ae2324b),
	.w4(32'hba372464),
	.w5(32'h3aa15cc8),
	.w6(32'h3aec7271),
	.w7(32'hbb94b978),
	.w8(32'hbb739604),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb21d7ba),
	.w1(32'h3bcef5fe),
	.w2(32'h3b9d20c0),
	.w3(32'hbb5ee0e0),
	.w4(32'h3a728592),
	.w5(32'h3ae92b8e),
	.w6(32'hbc19f5c5),
	.w7(32'hbb2803e0),
	.w8(32'hbb85dd79),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0390fe),
	.w1(32'h3981dff7),
	.w2(32'h3a0c3c72),
	.w3(32'hba0341c7),
	.w4(32'hba5d1796),
	.w5(32'hbb50a782),
	.w6(32'hbb247285),
	.w7(32'h3ace5f1f),
	.w8(32'h3b200a13),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afafc8f),
	.w1(32'hbbafd704),
	.w2(32'h3b01a662),
	.w3(32'h3af178ec),
	.w4(32'hbb5500fa),
	.w5(32'h3c347653),
	.w6(32'h3a00a31a),
	.w7(32'hbb294e42),
	.w8(32'h3a80d62d),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ada25a1),
	.w1(32'hbbe1176b),
	.w2(32'hbbfba79f),
	.w3(32'hbc084ce6),
	.w4(32'h3aada0bc),
	.w5(32'hbb1c3134),
	.w6(32'hbc433972),
	.w7(32'hbb882abe),
	.w8(32'hbb93270c),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb847f59b),
	.w1(32'hbbe0402d),
	.w2(32'hbb7154b4),
	.w3(32'h3b9f901f),
	.w4(32'h3bd240c1),
	.w5(32'h3b8524e2),
	.w6(32'hba3b4edd),
	.w7(32'h3aa08bb3),
	.w8(32'h3bf806a5),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb991d3d),
	.w1(32'hba9893c5),
	.w2(32'h3b4347f4),
	.w3(32'h3bd2f91f),
	.w4(32'h3b549cfc),
	.w5(32'hba6dc7ed),
	.w6(32'hb8e3d8d8),
	.w7(32'hbb31f229),
	.w8(32'h3887c4cb),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b49c7f8),
	.w1(32'hbb5fd0e4),
	.w2(32'h3b29b38e),
	.w3(32'hbbc1b899),
	.w4(32'h3b902a69),
	.w5(32'h3aca1dc6),
	.w6(32'hbb113605),
	.w7(32'h3a1c7b92),
	.w8(32'h3ba203a8),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa63a56),
	.w1(32'hbc027f8a),
	.w2(32'h3aa31980),
	.w3(32'h3b9ad996),
	.w4(32'hbc71c76b),
	.w5(32'hbc6d0529),
	.w6(32'h3bf3564a),
	.w7(32'hbc2f6a84),
	.w8(32'hbbf08334),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1b75b8),
	.w1(32'hbb0d2df2),
	.w2(32'h3b879b6a),
	.w3(32'hbbd78502),
	.w4(32'hbb54ea4a),
	.w5(32'h3bb72b9b),
	.w6(32'h3a47959b),
	.w7(32'hbb6bae23),
	.w8(32'h3b3b8d59),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c28de13),
	.w1(32'h3bb34a5c),
	.w2(32'h3c56b9ce),
	.w3(32'hbb84a746),
	.w4(32'h3bd79b2e),
	.w5(32'h3c964e39),
	.w6(32'hbb782b61),
	.w7(32'hbbf3928c),
	.w8(32'h3bcb1191),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b690002),
	.w1(32'h3b4a90fd),
	.w2(32'h3c03da1d),
	.w3(32'h3b71193c),
	.w4(32'h3a907737),
	.w5(32'h3c66c57d),
	.w6(32'h3b3f52f8),
	.w7(32'hbaf35ed9),
	.w8(32'h3c1bf134),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc35e59b),
	.w1(32'h3c0464e2),
	.w2(32'h3b682842),
	.w3(32'hbbb93aae),
	.w4(32'h3b90ead9),
	.w5(32'h3bbcbb84),
	.w6(32'h3bec80c6),
	.w7(32'h3ba6d159),
	.w8(32'h3c43ce74),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4fa063),
	.w1(32'hbbf59899),
	.w2(32'hbad1f0a9),
	.w3(32'h3a6de5f1),
	.w4(32'hbc15d41c),
	.w5(32'hbb87f319),
	.w6(32'h3b9b16bb),
	.w7(32'hbbc6b390),
	.w8(32'hbb8c197f),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2a3440),
	.w1(32'h3bd5845f),
	.w2(32'h3ac93b64),
	.w3(32'hbbd4e36d),
	.w4(32'h3be22321),
	.w5(32'h3c7198fc),
	.w6(32'hbb436eda),
	.w7(32'hbb21d0cd),
	.w8(32'h3c4134c3),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5d1638),
	.w1(32'h3add16f1),
	.w2(32'hba653c64),
	.w3(32'h3c255c6c),
	.w4(32'h3ba17d0c),
	.w5(32'hb998f28a),
	.w6(32'hb7ad7b99),
	.w7(32'h39d9b3c3),
	.w8(32'h3ab91390),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8044a4),
	.w1(32'h3acbda4f),
	.w2(32'h3c161981),
	.w3(32'hbb9fcbbf),
	.w4(32'hb9ab5656),
	.w5(32'h3bb409a6),
	.w6(32'hbb36ccd5),
	.w7(32'h3b92f86b),
	.w8(32'h3c1d09f7),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8d274e),
	.w1(32'hbc3a90c8),
	.w2(32'hbc5971b7),
	.w3(32'hbac921f0),
	.w4(32'hba96e7f6),
	.w5(32'hbc98f0cb),
	.w6(32'hbab6bddc),
	.w7(32'h3bb95e34),
	.w8(32'h3bc56958),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8aa1e2),
	.w1(32'hbb6c5fef),
	.w2(32'h3b1c8fbd),
	.w3(32'hb90db0f4),
	.w4(32'h3bdd8103),
	.w5(32'hba9e82d1),
	.w6(32'hbbd8cd23),
	.w7(32'h3b9eeceb),
	.w8(32'h3bda22a6),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3dad00),
	.w1(32'h3a581a1b),
	.w2(32'h3c4b691b),
	.w3(32'h38b1afee),
	.w4(32'h3cc1840e),
	.w5(32'h3d116942),
	.w6(32'h3ad9d4e3),
	.w7(32'h3c57b33a),
	.w8(32'h3cb9329a),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbba797),
	.w1(32'hbb45da92),
	.w2(32'hbbc75dad),
	.w3(32'h3ca896f9),
	.w4(32'h3bf5fd4f),
	.w5(32'h3c90505a),
	.w6(32'h3c433353),
	.w7(32'hb9350068),
	.w8(32'h3aea688d),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1028d7),
	.w1(32'hbbc728b1),
	.w2(32'hbac20245),
	.w3(32'hbb241e9c),
	.w4(32'h3b7d2b20),
	.w5(32'hbb8f8b30),
	.w6(32'hbbbf005c),
	.w7(32'h3ba9b2bd),
	.w8(32'h3c0cfddf),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2df9f5),
	.w1(32'h38f4ba05),
	.w2(32'h3b87f6b3),
	.w3(32'h3a3a623b),
	.w4(32'h39c4c14b),
	.w5(32'hbb9aff45),
	.w6(32'hbb0f6650),
	.w7(32'hbacd5fb4),
	.w8(32'hbb42ee57),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc5f93e),
	.w1(32'h3bfcd4b5),
	.w2(32'hbc06175a),
	.w3(32'hbb3d0004),
	.w4(32'h3b1207c3),
	.w5(32'hbc0dd309),
	.w6(32'hbb06e5fd),
	.w7(32'h3b820ed3),
	.w8(32'h3ac0092e),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb23e68),
	.w1(32'h3a0750a6),
	.w2(32'h3b8e4754),
	.w3(32'h399169e7),
	.w4(32'hba6fa0db),
	.w5(32'h3b19f907),
	.w6(32'h3c18b11e),
	.w7(32'h3ac4f6c5),
	.w8(32'hbb1e1c18),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b25cc23),
	.w1(32'hbb39e400),
	.w2(32'h3aca0899),
	.w3(32'hbb0b56c6),
	.w4(32'hbb6336ae),
	.w5(32'h3a8856bc),
	.w6(32'h3b0e1480),
	.w7(32'hba4fac14),
	.w8(32'hbba971ee),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1c0feb),
	.w1(32'h3bcfc3f4),
	.w2(32'h3c0bfbc3),
	.w3(32'h3bc44b30),
	.w4(32'hb9fdd221),
	.w5(32'hbb0814b1),
	.w6(32'hbaec8266),
	.w7(32'h3bcf9d81),
	.w8(32'h3ab3120b),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c22e03c),
	.w1(32'hbb19f810),
	.w2(32'h3bd0f357),
	.w3(32'h3b2cde1b),
	.w4(32'hbb2f80d1),
	.w5(32'hbb5fa3f6),
	.w6(32'h3a5a3d0b),
	.w7(32'hbabc5b98),
	.w8(32'h3bd14262),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1bee1e),
	.w1(32'hbbfb1699),
	.w2(32'hbb81fc74),
	.w3(32'h3bbfe45a),
	.w4(32'h3a3c9114),
	.w5(32'hbb8ef838),
	.w6(32'h3bbcab44),
	.w7(32'hbabe8cc7),
	.w8(32'h3a0bc41f),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba924bc3),
	.w1(32'hbae9eb07),
	.w2(32'h3bd24cc8),
	.w3(32'hbbdfd611),
	.w4(32'hbc40563a),
	.w5(32'h3c162988),
	.w6(32'hbbba16c1),
	.w7(32'hba4043c0),
	.w8(32'hbc4ed990),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaca4d29),
	.w1(32'h3b3beed4),
	.w2(32'h3b12c75e),
	.w3(32'h3bd6ace6),
	.w4(32'h3af2b55b),
	.w5(32'hbb8c2143),
	.w6(32'h3b11d80c),
	.w7(32'h3b31af5c),
	.w8(32'h3b42055f),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6f84ee),
	.w1(32'hbb47ca5e),
	.w2(32'h3b6a640b),
	.w3(32'hbbcb819a),
	.w4(32'h3b1b1133),
	.w5(32'h3b6f86d8),
	.w6(32'hbb8c4589),
	.w7(32'h37763105),
	.w8(32'hbc1cbab7),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb043946),
	.w1(32'hbb1feea9),
	.w2(32'h3ba92989),
	.w3(32'hbb8aca6c),
	.w4(32'h3a2caecb),
	.w5(32'hba2b48ca),
	.w6(32'hbc1ef976),
	.w7(32'hbb57c4e3),
	.w8(32'hbc12cead),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb220b5a),
	.w1(32'h3c0f5a6a),
	.w2(32'h3c07cd92),
	.w3(32'hbc0fa228),
	.w4(32'h3c09403a),
	.w5(32'hbaafcf0a),
	.w6(32'hbb3e2a2f),
	.w7(32'h3c83789c),
	.w8(32'h3c0031da),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c340b0c),
	.w1(32'hbb5cbce3),
	.w2(32'hbc203efc),
	.w3(32'h3b0f1bf5),
	.w4(32'hbc56870f),
	.w5(32'hbc5a8806),
	.w6(32'h3c19fcf0),
	.w7(32'hbc5805ab),
	.w8(32'hbc429b2a),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4a86a7),
	.w1(32'hb969dab3),
	.w2(32'h3b91cadc),
	.w3(32'hbc13398f),
	.w4(32'hbbb8e000),
	.w5(32'h3b27c65b),
	.w6(32'hba891cff),
	.w7(32'hbb2b7b0b),
	.w8(32'h3bee767f),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb701c3),
	.w1(32'hbb1e316a),
	.w2(32'hbaf46417),
	.w3(32'h3b1f228a),
	.w4(32'hbbf22e2d),
	.w5(32'hbabc7c72),
	.w6(32'hbb5836b3),
	.w7(32'h3b608f10),
	.w8(32'h3c1a1ad5),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb92dde1),
	.w1(32'hb7facaca),
	.w2(32'h3abac50a),
	.w3(32'hbc097fc7),
	.w4(32'h3b8ef1f1),
	.w5(32'h3b819c56),
	.w6(32'h3c215718),
	.w7(32'h3c207b3d),
	.w8(32'h3bb92cf0),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0a2bfe),
	.w1(32'hbaafd467),
	.w2(32'hbb7a8eb0),
	.w3(32'h3bcb9358),
	.w4(32'hbab6edb1),
	.w5(32'hbc036de3),
	.w6(32'h3abcb330),
	.w7(32'h3a92f78d),
	.w8(32'h3b4ce6d8),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac94807),
	.w1(32'h3b2ed790),
	.w2(32'hbaf901a6),
	.w3(32'h3aed881e),
	.w4(32'h3a171f87),
	.w5(32'hbc16083a),
	.w6(32'h3bffaaba),
	.w7(32'h38acbf03),
	.w8(32'h3b1da327),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb0726b),
	.w1(32'h3a91c8d1),
	.w2(32'h3be6cddd),
	.w3(32'hba1b3642),
	.w4(32'hbc1850cc),
	.w5(32'hbb5d8702),
	.w6(32'h3969a4a8),
	.w7(32'hbbe45403),
	.w8(32'h3a4d16f1),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8f28fb),
	.w1(32'h3b4c40ce),
	.w2(32'hbaeea452),
	.w3(32'h39789d97),
	.w4(32'hb9412cdd),
	.w5(32'h3b60ea8e),
	.w6(32'hbc154233),
	.w7(32'h3857ca94),
	.w8(32'h3c151cd3),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a627712),
	.w1(32'hb63a3f9c),
	.w2(32'h3b5c61f2),
	.w3(32'hbb4051d6),
	.w4(32'h3c8c378f),
	.w5(32'h3cc82a83),
	.w6(32'h3b548f6b),
	.w7(32'h3c9554e1),
	.w8(32'h3cf4bd9d),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6cbf20),
	.w1(32'h3b4b58aa),
	.w2(32'h3afb8c7b),
	.w3(32'h3c0ee0fa),
	.w4(32'h3c8acff9),
	.w5(32'h3c78574c),
	.w6(32'h3c402b70),
	.w7(32'h3bf5c692),
	.w8(32'h3a85877a),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0d103d),
	.w1(32'h3b070281),
	.w2(32'hbb9072a4),
	.w3(32'h3c5ba019),
	.w4(32'h3b5d4904),
	.w5(32'hbc857b51),
	.w6(32'hbb380582),
	.w7(32'h3c477355),
	.w8(32'h3c50c7d8),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb31cf9b),
	.w1(32'hbbc0f7fe),
	.w2(32'hba9e83a5),
	.w3(32'hba856d2c),
	.w4(32'hb9d2db40),
	.w5(32'hbb858ce9),
	.w6(32'hbb05661c),
	.w7(32'h3b0565e1),
	.w8(32'hbb2abb9d),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa12eb5),
	.w1(32'h3abac771),
	.w2(32'h39e6b714),
	.w3(32'hbac68915),
	.w4(32'hbb1c2786),
	.w5(32'h3c251aeb),
	.w6(32'hbbb5c8b5),
	.w7(32'hbbb89ccb),
	.w8(32'hba6e3e2d),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdb428e),
	.w1(32'hbb1f8418),
	.w2(32'hbb6caacc),
	.w3(32'hbc039bf1),
	.w4(32'hb950f3f2),
	.w5(32'h3b2690bd),
	.w6(32'hbb9c7b52),
	.w7(32'h3b5a81d5),
	.w8(32'hba4cc7b9),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba58b35),
	.w1(32'h3b58abdc),
	.w2(32'h3c1050d0),
	.w3(32'hbaa69bb9),
	.w4(32'h3b5dfa00),
	.w5(32'h3b2b743d),
	.w6(32'h39fc664b),
	.w7(32'h38a19a05),
	.w8(32'h3a8193a2),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aac48b8),
	.w1(32'hbac09d7c),
	.w2(32'hbb0baeb2),
	.w3(32'h3bdc0db9),
	.w4(32'hbb472108),
	.w5(32'hbb8ecd8e),
	.w6(32'h3b541db8),
	.w7(32'h3bde344f),
	.w8(32'h3b58143f),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5f6523),
	.w1(32'hbc2dafc0),
	.w2(32'hbbb80999),
	.w3(32'hbb2b5883),
	.w4(32'hbb962cd1),
	.w5(32'hbc3244db),
	.w6(32'h3ad9f498),
	.w7(32'h3bd7ef99),
	.w8(32'h3b4b318d),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba89e2e1),
	.w1(32'hb858f16a),
	.w2(32'hbbf2a9e4),
	.w3(32'hbb5ff9ea),
	.w4(32'hbb1cd422),
	.w5(32'hbb3f83e6),
	.w6(32'h3b89524d),
	.w7(32'hbaaf3673),
	.w8(32'h3b1b47e8),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba0839e),
	.w1(32'h3b505b22),
	.w2(32'hbb3a36b0),
	.w3(32'hbbe832b8),
	.w4(32'hb9fce2c5),
	.w5(32'hbb94d70f),
	.w6(32'hb9fcf0b1),
	.w7(32'h3b969af8),
	.w8(32'h3c05f127),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba68c241),
	.w1(32'h3b6836cd),
	.w2(32'h3c1716ef),
	.w3(32'hbb6853f1),
	.w4(32'hbaea5084),
	.w5(32'h3bad9e80),
	.w6(32'h3bdf30ed),
	.w7(32'hba92aaa7),
	.w8(32'h3b149d34),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b89483e),
	.w1(32'h3b1fb632),
	.w2(32'h3c0e2196),
	.w3(32'h3b706fc7),
	.w4(32'h3b830f13),
	.w5(32'h3c11d58c),
	.w6(32'h3b74df02),
	.w7(32'h3bea375a),
	.w8(32'h3bc3e7c9),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a081794),
	.w1(32'hbb2cb79b),
	.w2(32'h3a4fdf6f),
	.w3(32'h3b53829e),
	.w4(32'hb79642d0),
	.w5(32'h3ab716aa),
	.w6(32'h3adc7238),
	.w7(32'h3be982c1),
	.w8(32'h3b1354e3),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0e0eb6),
	.w1(32'h3aa2ecdd),
	.w2(32'h3c64e523),
	.w3(32'h3b4da91e),
	.w4(32'hbab44c33),
	.w5(32'h3a1f54e4),
	.w6(32'hb9b94043),
	.w7(32'hbbcfc02e),
	.w8(32'hbb2c3395),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a4ed2eb),
	.w1(32'h3b408640),
	.w2(32'h3abeb369),
	.w3(32'hbbcc14c3),
	.w4(32'h3adddf31),
	.w5(32'hbbbb178d),
	.w6(32'hbb2cf037),
	.w7(32'hbb0351d5),
	.w8(32'h37edcebd),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4e3fb7),
	.w1(32'h3b021627),
	.w2(32'hbb195e77),
	.w3(32'h3a5bd136),
	.w4(32'h3bd9b890),
	.w5(32'hbbc27dc3),
	.w6(32'hbb64581c),
	.w7(32'h3ad639bb),
	.w8(32'h3bb340d0),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb6f2aa),
	.w1(32'hbbc5dd06),
	.w2(32'hbbbb2325),
	.w3(32'h39bd2b08),
	.w4(32'h3af700f8),
	.w5(32'hba61353a),
	.w6(32'hbbe9b169),
	.w7(32'h3abfe170),
	.w8(32'h3c45ed08),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb54b3f3),
	.w1(32'hbb487818),
	.w2(32'hb9c8dbf6),
	.w3(32'h3bb2d39f),
	.w4(32'h3b6969c0),
	.w5(32'hbbee5503),
	.w6(32'hbb828cc5),
	.w7(32'hba5eeac6),
	.w8(32'h3bd5762b),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5a5d7a),
	.w1(32'h3ba0746d),
	.w2(32'h3c0614e4),
	.w3(32'h3b232bfd),
	.w4(32'h3c02b064),
	.w5(32'h3c95edfe),
	.w6(32'h3ba901c9),
	.w7(32'h3abbbc78),
	.w8(32'h3b39be19),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4e808e),
	.w1(32'hb8c6171f),
	.w2(32'h3ab2177e),
	.w3(32'h3bb13668),
	.w4(32'hbbaa80a4),
	.w5(32'hbc52bb39),
	.w6(32'hbb5d908e),
	.w7(32'h3bcc9d6a),
	.w8(32'h3b549260),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a790267),
	.w1(32'h3aa86f3f),
	.w2(32'hbb711bc2),
	.w3(32'hbb086284),
	.w4(32'hbb67b4bd),
	.w5(32'hbc16f847),
	.w6(32'hbb6c2f6a),
	.w7(32'h3b8d087a),
	.w8(32'h3ad0d4bb),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc39484f),
	.w1(32'hbb627e58),
	.w2(32'hbc0fed98),
	.w3(32'hbc2b0f82),
	.w4(32'h3a5a5b01),
	.w5(32'hb9360ea7),
	.w6(32'hbb43055e),
	.w7(32'h3c777396),
	.w8(32'h3c54aa91),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba81901a),
	.w1(32'h3bb89dd9),
	.w2(32'h3bfa7d20),
	.w3(32'hba3383b4),
	.w4(32'h3b56e79b),
	.w5(32'h3b86be2a),
	.w6(32'h3beba2fa),
	.w7(32'h3c0d61f8),
	.w8(32'h3c28ea62),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8ba88e),
	.w1(32'h3b67f3ba),
	.w2(32'h3c436b20),
	.w3(32'h3ad9d851),
	.w4(32'hba9da4e6),
	.w5(32'h3c588c73),
	.w6(32'h3befb6c1),
	.w7(32'hbc08a70e),
	.w8(32'h3b812ed7),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3f0256),
	.w1(32'hbaa57a46),
	.w2(32'h3bb36ebb),
	.w3(32'h3c247a90),
	.w4(32'h3a57c2b8),
	.w5(32'h3c6ecd2f),
	.w6(32'h3be16044),
	.w7(32'hbc088361),
	.w8(32'h3c3a3664),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6ff255),
	.w1(32'h3ba49a63),
	.w2(32'h3b755332),
	.w3(32'h3b5a1a02),
	.w4(32'h3b936320),
	.w5(32'h3b9064e1),
	.w6(32'h3b0d1143),
	.w7(32'h3c84dc73),
	.w8(32'hba9e5eaa),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c633d4e),
	.w1(32'h3c8f55be),
	.w2(32'h3d20ac96),
	.w3(32'h3c5b465e),
	.w4(32'h3bb9e131),
	.w5(32'h3caadf7e),
	.w6(32'h3c8ef19d),
	.w7(32'hbb3e8eb6),
	.w8(32'h3c037061),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5bf61c),
	.w1(32'h3b836a19),
	.w2(32'h3a1423e2),
	.w3(32'h3c9bdc4b),
	.w4(32'h3bacbcc8),
	.w5(32'hbb9af472),
	.w6(32'h3a9298b9),
	.w7(32'h3c0a6e94),
	.w8(32'h3cbd7720),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac80b85),
	.w1(32'hbb4fb8bf),
	.w2(32'hbb9daf6a),
	.w3(32'h3b038324),
	.w4(32'h3b9919c8),
	.w5(32'hb88748e1),
	.w6(32'h3c0aa69a),
	.w7(32'h3c0b2f3e),
	.w8(32'h3c2e5d7a),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb236ed3),
	.w1(32'hba9a8280),
	.w2(32'h3b3a0da3),
	.w3(32'h39a5e9d4),
	.w4(32'hbb6de9d4),
	.w5(32'hbc013360),
	.w6(32'h3b36cc51),
	.w7(32'hbaf2c61d),
	.w8(32'hbb80f016),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b434102),
	.w1(32'hbb595f3c),
	.w2(32'h3b1cd301),
	.w3(32'hbb7c23a6),
	.w4(32'h3c390661),
	.w5(32'h3babbcb8),
	.w6(32'h3af895df),
	.w7(32'hb96a2195),
	.w8(32'h3c29df9d),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2caf4e),
	.w1(32'h3a23bfd0),
	.w2(32'h3ac09446),
	.w3(32'h3c100d86),
	.w4(32'h3bf8dc69),
	.w5(32'h3c303800),
	.w6(32'h3b2e4110),
	.w7(32'hb9e2698a),
	.w8(32'h3b615e08),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9cd2a6),
	.w1(32'hbaf35b2a),
	.w2(32'hbb8c25b0),
	.w3(32'h3c17d089),
	.w4(32'hbb7aa13c),
	.w5(32'hbb9c81cb),
	.w6(32'h3b8c2615),
	.w7(32'h3b075139),
	.w8(32'h3a8ea3dc),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb61da33),
	.w1(32'hbb4444e8),
	.w2(32'hbbb2eae0),
	.w3(32'hbc029f94),
	.w4(32'hba92dc46),
	.w5(32'hbac13704),
	.w6(32'hbb9074a8),
	.w7(32'hbb9e85ca),
	.w8(32'h3b96bc57),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba7d4d7),
	.w1(32'h3b283841),
	.w2(32'hbba2eb69),
	.w3(32'hbbf9832c),
	.w4(32'h3bc50cf2),
	.w5(32'hbbbfc345),
	.w6(32'hbc895b46),
	.w7(32'hbc89e264),
	.w8(32'h3c803ec5),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb733aa2),
	.w1(32'h3885f155),
	.w2(32'h3b59d4be),
	.w3(32'hbab87196),
	.w4(32'hbbcce67c),
	.w5(32'hbb519369),
	.w6(32'h3bcfd57f),
	.w7(32'hbc054e4d),
	.w8(32'hbb9cfa57),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc783691),
	.w1(32'hbc96e240),
	.w2(32'hba6a1387),
	.w3(32'hbc3a62dd),
	.w4(32'hbc95221c),
	.w5(32'hbc3c85b8),
	.w6(32'hbbd68d80),
	.w7(32'hbbec416e),
	.w8(32'hbc7a71aa),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae46dc7),
	.w1(32'h3a782081),
	.w2(32'h3c1af7d2),
	.w3(32'hbbf91a1a),
	.w4(32'hb9f5e527),
	.w5(32'h3a94d06c),
	.w6(32'hbc74727f),
	.w7(32'h3aa7d37e),
	.w8(32'h3c2ba0ea),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a02e079),
	.w1(32'hbc1f6c98),
	.w2(32'hbbd53986),
	.w3(32'hb9d4ee81),
	.w4(32'hbbba3763),
	.w5(32'h3c3e3b6b),
	.w6(32'h3b526e0a),
	.w7(32'h3b84e15d),
	.w8(32'h3bf318dd),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b091856),
	.w1(32'hbb23c2d7),
	.w2(32'hbc061747),
	.w3(32'h3c141362),
	.w4(32'hbab95b87),
	.w5(32'hbb154408),
	.w6(32'h3c352fe7),
	.w7(32'h3ab0f493),
	.w8(32'hbbfd840f),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc28513),
	.w1(32'hba12736e),
	.w2(32'h3a90689f),
	.w3(32'hbbb6cc32),
	.w4(32'h3a8746c8),
	.w5(32'h3b110f3b),
	.w6(32'hba414fbc),
	.w7(32'hbb92981e),
	.w8(32'hbc0c4810),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af8bd5a),
	.w1(32'h3b9160a7),
	.w2(32'hbaa2914b),
	.w3(32'hba14854e),
	.w4(32'hbaaf1ce7),
	.w5(32'h3cd86a67),
	.w6(32'hbb9b147a),
	.w7(32'h3b572a2f),
	.w8(32'h3c4930dd),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3bcdc1),
	.w1(32'hbb5261d9),
	.w2(32'hbbea6a17),
	.w3(32'h3c542280),
	.w4(32'h3abfcfb2),
	.w5(32'h3be2f5ca),
	.w6(32'h3c43fb70),
	.w7(32'h3bbfaf91),
	.w8(32'h3bd39634),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a450fe1),
	.w1(32'hbb9f8364),
	.w2(32'hbc1df3f8),
	.w3(32'h3be56ae3),
	.w4(32'hbb64580b),
	.w5(32'hbc386808),
	.w6(32'h3bc8e7c9),
	.w7(32'hbbfa42c7),
	.w8(32'hbbca29de),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba048eaa),
	.w1(32'hbab30678),
	.w2(32'h3a9b71b2),
	.w3(32'hbb36ca97),
	.w4(32'hbc55abae),
	.w5(32'h3ac2fbfd),
	.w6(32'h3b48b622),
	.w7(32'h39932dde),
	.w8(32'hbaac7afa),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c566986),
	.w1(32'hbbfabb91),
	.w2(32'hbc2b7176),
	.w3(32'h3b2964d0),
	.w4(32'hbb41280b),
	.w5(32'hbbb43a87),
	.w6(32'h3b9b3a98),
	.w7(32'hbb6bf566),
	.w8(32'h3a958d89),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac62fb8),
	.w1(32'h3b18e49d),
	.w2(32'hbbbb2e8b),
	.w3(32'h3be265c7),
	.w4(32'h3b230ae9),
	.w5(32'h3bd564b4),
	.w6(32'h39a0e72c),
	.w7(32'hbc52eb3c),
	.w8(32'h3c52074a),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2713e1),
	.w1(32'h3caec9f8),
	.w2(32'h3c7e3652),
	.w3(32'hbca9f9d9),
	.w4(32'hbb24bdb2),
	.w5(32'hbc950d57),
	.w6(32'hbbdbf296),
	.w7(32'hbc61d179),
	.w8(32'hbc571ff2),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c13a193),
	.w1(32'hb91e8726),
	.w2(32'hbacc20e1),
	.w3(32'hba72d67d),
	.w4(32'hbb76ce0f),
	.w5(32'hb949ddc2),
	.w6(32'hbb9badec),
	.w7(32'hbbd40c69),
	.w8(32'h3abcb3ff),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbca02bb),
	.w1(32'hbb55b810),
	.w2(32'hbbbab580),
	.w3(32'hba9dc277),
	.w4(32'h3ba0fd4b),
	.w5(32'h3bac5e9f),
	.w6(32'hb95ade82),
	.w7(32'hbae1888a),
	.w8(32'h3a72dde3),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe735f9),
	.w1(32'hbbc242aa),
	.w2(32'h3b658cbb),
	.w3(32'hbabed788),
	.w4(32'hbb82a193),
	.w5(32'h3c92624d),
	.w6(32'hbae2cec0),
	.w7(32'hbc382573),
	.w8(32'h3c121584),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c17396a),
	.w1(32'hbbf71620),
	.w2(32'hbbc8ab4d),
	.w3(32'h3c0607d9),
	.w4(32'hbbbd63ed),
	.w5(32'h3b7e17b6),
	.w6(32'hb94af1c3),
	.w7(32'h3b91f386),
	.w8(32'h3c046b81),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39ad9585),
	.w1(32'h3ba93047),
	.w2(32'h3c22ad84),
	.w3(32'h3b96e673),
	.w4(32'h3bb43c63),
	.w5(32'h3be9e013),
	.w6(32'h3b3cd164),
	.w7(32'h3c62cfee),
	.w8(32'hbb26e80a),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baea1f2),
	.w1(32'h3bb4800d),
	.w2(32'h3b72808d),
	.w3(32'hbb94059b),
	.w4(32'h3b9f4830),
	.w5(32'h3c686218),
	.w6(32'hbbc1a0cf),
	.w7(32'hbc02697d),
	.w8(32'h3bf53d70),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb90c138),
	.w1(32'hbba25bd2),
	.w2(32'h3a9116a9),
	.w3(32'h3b5881e1),
	.w4(32'h3c26aab3),
	.w5(32'h3cb1ca0c),
	.w6(32'h3bade0f5),
	.w7(32'hbba2b1a4),
	.w8(32'hbb67bb5d),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb2cb50),
	.w1(32'hbc1979ef),
	.w2(32'hbc480cc0),
	.w3(32'h3b7fcecb),
	.w4(32'hbc018cd3),
	.w5(32'hbb62818a),
	.w6(32'hbb17038a),
	.w7(32'h3b4d3626),
	.w8(32'h3c8e50bc),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb90b813),
	.w1(32'hbb85087b),
	.w2(32'h3a3891ed),
	.w3(32'hbb9a7747),
	.w4(32'hb9f7c001),
	.w5(32'hbb9525a1),
	.w6(32'h3bd94a28),
	.w7(32'hbc301724),
	.w8(32'hbbfc7f92),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc146056),
	.w1(32'hbb8578d0),
	.w2(32'h3c610abe),
	.w3(32'hbbb25082),
	.w4(32'hbbcff62f),
	.w5(32'h3b98706b),
	.w6(32'hbbf7fca7),
	.w7(32'hbbe84ba4),
	.w8(32'hba6b5daf),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba2abb2),
	.w1(32'h3c01cdd2),
	.w2(32'h3c4a953e),
	.w3(32'hbc2cad7e),
	.w4(32'h3c956bc6),
	.w5(32'h3cc50de8),
	.w6(32'hbb7d11ed),
	.w7(32'h3b811f37),
	.w8(32'h3b974de5),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c54169f),
	.w1(32'hba95f001),
	.w2(32'hbc1d4624),
	.w3(32'h3caf7ced),
	.w4(32'hbba4bfaf),
	.w5(32'hbbdb6a4d),
	.w6(32'h3c1e8081),
	.w7(32'hbbe93cb4),
	.w8(32'hbc221a6e),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4e3c85),
	.w1(32'hbb662766),
	.w2(32'hbc1a84f4),
	.w3(32'h3a53450c),
	.w4(32'h3ace5d1c),
	.w5(32'hbc6a4c03),
	.w6(32'hbbc14efa),
	.w7(32'hbba171af),
	.w8(32'hbc225f94),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb59ca80),
	.w1(32'h3b9005a0),
	.w2(32'hbbabaea2),
	.w3(32'hba3d7d5d),
	.w4(32'h3c950ccc),
	.w5(32'h3cbd1592),
	.w6(32'hbbacb9ba),
	.w7(32'h3c9ceef7),
	.w8(32'h3ce55d48),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa8e032),
	.w1(32'h3a6a615c),
	.w2(32'hbc59f849),
	.w3(32'h3c442fd3),
	.w4(32'hbc498380),
	.w5(32'h3aa16613),
	.w6(32'h3ca5353a),
	.w7(32'hbbc1ab61),
	.w8(32'hbbaed9e4),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc663139),
	.w1(32'hbabe2804),
	.w2(32'h3bf6b0f2),
	.w3(32'hbc2d10be),
	.w4(32'hbb6bacf2),
	.w5(32'h3bab5164),
	.w6(32'h3a2d1626),
	.w7(32'hbb73f5df),
	.w8(32'h3a2fa916),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c042aaa),
	.w1(32'hbb8fc811),
	.w2(32'hbabd2ecc),
	.w3(32'h3bad458f),
	.w4(32'hbac9deb4),
	.w5(32'hbbf734c7),
	.w6(32'h3a7da231),
	.w7(32'hbb4ecae9),
	.w8(32'hbc0a9853),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0ce78e),
	.w1(32'hbc25f8b8),
	.w2(32'hbc11c5d6),
	.w3(32'hbbe38216),
	.w4(32'hbb843288),
	.w5(32'hbb9e2b6c),
	.w6(32'hbc2fb7a1),
	.w7(32'h3bcbdf29),
	.w8(32'h3bd4f138),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1b8393),
	.w1(32'h3b89c232),
	.w2(32'h3bf7103a),
	.w3(32'hba719af3),
	.w4(32'hbc7ffb84),
	.w5(32'hbc40834e),
	.w6(32'hbb1344ae),
	.w7(32'hbba576eb),
	.w8(32'hbbe245bf),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c54503b),
	.w1(32'h3b014b86),
	.w2(32'hbad3b64a),
	.w3(32'hbc6399d9),
	.w4(32'hbac7a746),
	.w5(32'h39d6feaf),
	.w6(32'hbb4ce008),
	.w7(32'h3a3028f5),
	.w8(32'h3c19304c),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9533a7),
	.w1(32'hbc0756dd),
	.w2(32'hbb7632aa),
	.w3(32'h3ba352ba),
	.w4(32'h3af73afe),
	.w5(32'hbb0d9c12),
	.w6(32'h3badd2f7),
	.w7(32'h3aaf91fd),
	.w8(32'hbbf4ddac),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc6f500),
	.w1(32'hbc7b1fd0),
	.w2(32'hbb2877e8),
	.w3(32'hbc059c9c),
	.w4(32'hbb9c92bc),
	.w5(32'h3c9bf391),
	.w6(32'hbc021f34),
	.w7(32'hbbd77e67),
	.w8(32'hbb371673),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395a3a2e),
	.w1(32'hbb7f98b3),
	.w2(32'hbb63ffd9),
	.w3(32'h3c0bf26f),
	.w4(32'h3abf41ae),
	.w5(32'h3b0298ec),
	.w6(32'h3b9ad905),
	.w7(32'hbb8d3d95),
	.w8(32'hb9071a8f),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb36d9d3),
	.w1(32'hbb963022),
	.w2(32'h3b359784),
	.w3(32'h3b8a51f4),
	.w4(32'h3c55fac5),
	.w5(32'h3c2b0ce2),
	.w6(32'h3bbd98fb),
	.w7(32'h3c34ab9a),
	.w8(32'h3bec44b8),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab56303),
	.w1(32'hbbd18ca4),
	.w2(32'hbb5071d7),
	.w3(32'hbb9e6e4e),
	.w4(32'hbc0834b8),
	.w5(32'hbb383337),
	.w6(32'h3aeaa8bc),
	.w7(32'h3ba67336),
	.w8(32'h3c28e9df),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3a8922),
	.w1(32'h3ba8d021),
	.w2(32'h3bad58f6),
	.w3(32'h3b756714),
	.w4(32'h3b877f7e),
	.w5(32'hba28c2fc),
	.w6(32'h3c07e6e2),
	.w7(32'hb9731810),
	.w8(32'hbb5b83ac),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba62d35e),
	.w1(32'hbbe875c6),
	.w2(32'h3c24de75),
	.w3(32'hbb8c095a),
	.w4(32'hbb8389bb),
	.w5(32'hb7f33f5f),
	.w6(32'hbbb9357b),
	.w7(32'hbb869506),
	.w8(32'hbc0f11ce),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c23f2ee),
	.w1(32'hbb4d07d7),
	.w2(32'h3921a77d),
	.w3(32'h3c15f681),
	.w4(32'hbbcf2c63),
	.w5(32'h3b703411),
	.w6(32'hbb86e359),
	.w7(32'hbc097590),
	.w8(32'hbb63507b),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aba2d85),
	.w1(32'hbbede911),
	.w2(32'hbc1837f3),
	.w3(32'h3b0474a8),
	.w4(32'h3bf152b4),
	.w5(32'h3c3de7e6),
	.w6(32'hbbc14aed),
	.w7(32'hb83bae19),
	.w8(32'h3be76769),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2a8241),
	.w1(32'h3ca286c2),
	.w2(32'h3cecded0),
	.w3(32'h39b91b02),
	.w4(32'h3c61cbb7),
	.w5(32'hba3caf04),
	.w6(32'h3bba0172),
	.w7(32'hbac9e36f),
	.w8(32'hbb3539af),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c049b88),
	.w1(32'h3b5e5a1b),
	.w2(32'h3c7c3f3e),
	.w3(32'h3c5925af),
	.w4(32'h3a6deef5),
	.w5(32'h3ba0fc6a),
	.w6(32'hba4bc5eb),
	.w7(32'h3ad6e057),
	.w8(32'h3a41b94c),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4b2015),
	.w1(32'hbb825456),
	.w2(32'h3ae3d0ee),
	.w3(32'h3bbe07ae),
	.w4(32'h3b11deab),
	.w5(32'h3aaa6de6),
	.w6(32'h3ba5499d),
	.w7(32'h3a9809fd),
	.w8(32'h391f2447),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b60c40c),
	.w1(32'hbb534934),
	.w2(32'hbb4bc9b5),
	.w3(32'h3bcd1560),
	.w4(32'h3b462d85),
	.w5(32'h3bf39097),
	.w6(32'hb9a48a41),
	.w7(32'hbb18fa5d),
	.w8(32'h399835d7),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe176a6),
	.w1(32'hb9aba642),
	.w2(32'hbb90d246),
	.w3(32'h396bdd7f),
	.w4(32'h37897715),
	.w5(32'hbc109971),
	.w6(32'h3ab30fed),
	.w7(32'hbaf6f2a6),
	.w8(32'hbbe17f92),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a533157),
	.w1(32'hbc1608b9),
	.w2(32'hbc32892d),
	.w3(32'hbb7765ef),
	.w4(32'hbbd9659b),
	.w5(32'hbb7265f3),
	.w6(32'h39a38a4b),
	.w7(32'hbbbf9ce8),
	.w8(32'h3ace7a0f),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf51d56),
	.w1(32'hbab5d18e),
	.w2(32'hbbd08c26),
	.w3(32'h39b3db93),
	.w4(32'hbb59fb89),
	.w5(32'hb8c1a6d9),
	.w6(32'h3bcd5a41),
	.w7(32'hbc0fb162),
	.w8(32'hbc0787e8),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb949935),
	.w1(32'hbb3c416d),
	.w2(32'h3a94a089),
	.w3(32'h3b74b015),
	.w4(32'hbaa17dc2),
	.w5(32'hbc08d753),
	.w6(32'h3b8accd8),
	.w7(32'h3b47fd2b),
	.w8(32'hbbacd2b6),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94233d2),
	.w1(32'h3ba334aa),
	.w2(32'hba18d3bb),
	.w3(32'hbb59e13d),
	.w4(32'h3b292b53),
	.w5(32'h3c82de6a),
	.w6(32'hbaf17eae),
	.w7(32'hba88e5b5),
	.w8(32'h3b865779),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaadd4f2),
	.w1(32'hbbf65e00),
	.w2(32'hbb63a063),
	.w3(32'h3b9d14ff),
	.w4(32'hba24e856),
	.w5(32'h3b94bb16),
	.w6(32'h371f8f3f),
	.w7(32'hba29f88c),
	.w8(32'h3a365b4c),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae47577),
	.w1(32'hbb6e7d4a),
	.w2(32'hbbcf299a),
	.w3(32'h3b1e96e2),
	.w4(32'hba8e7422),
	.w5(32'hbb803bdb),
	.w6(32'hbb30653f),
	.w7(32'h3ab4679a),
	.w8(32'h3adbd92b),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7ae356),
	.w1(32'h3af1954c),
	.w2(32'hbb503aad),
	.w3(32'hbafe25d3),
	.w4(32'hbc33ff18),
	.w5(32'hbc41c9ab),
	.w6(32'h3b7c01a3),
	.w7(32'hbc5a9fca),
	.w8(32'hbc94652c),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd24183),
	.w1(32'hbb05e97b),
	.w2(32'h3ac1d964),
	.w3(32'hba5513c7),
	.w4(32'h3b6bf3d4),
	.w5(32'h3b976593),
	.w6(32'hbc6f3239),
	.w7(32'h3ba37cd4),
	.w8(32'h3c0fbc38),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b11bad8),
	.w1(32'h3bdba767),
	.w2(32'h3bf9c691),
	.w3(32'h3bab77ed),
	.w4(32'h3ac74407),
	.w5(32'hbb4282c3),
	.w6(32'hb95ee717),
	.w7(32'h3b4b65ea),
	.w8(32'hbb9cf652),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8e18ab),
	.w1(32'hbc179763),
	.w2(32'hbbabdb24),
	.w3(32'h3c777acb),
	.w4(32'hbc0b38ca),
	.w5(32'h3bd490c1),
	.w6(32'hbb1cb455),
	.w7(32'h3c1a4be3),
	.w8(32'h3c3b20c8),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab74e56),
	.w1(32'hbbdbbb42),
	.w2(32'h3b1cde9f),
	.w3(32'h3c2ee58b),
	.w4(32'h3c8a5832),
	.w5(32'h3d00ce58),
	.w6(32'h3c67c88f),
	.w7(32'h3c513147),
	.w8(32'h3c6587b4),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb996da56),
	.w1(32'h3c00f8b4),
	.w2(32'h3c260cdc),
	.w3(32'h3c340fb4),
	.w4(32'hbbce2afb),
	.w5(32'hb9c306ff),
	.w6(32'hbac1912a),
	.w7(32'h3bb75c28),
	.w8(32'h3c4c80f6),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c425e08),
	.w1(32'hbbe3076a),
	.w2(32'h3c30b874),
	.w3(32'h3b9ffe3a),
	.w4(32'hb90d8e36),
	.w5(32'h3cc84830),
	.w6(32'h3c90cfed),
	.w7(32'h3c13f56d),
	.w8(32'h3c871704),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule