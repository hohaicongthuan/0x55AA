module layer_10_featuremap_321(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac95644),
	.w1(32'hbabd868c),
	.w2(32'hb9835ba9),
	.w3(32'h39da01ac),
	.w4(32'h3942704c),
	.w5(32'hba8c1380),
	.w6(32'h399bad07),
	.w7(32'hb8fb16d9),
	.w8(32'hbb0af3cc),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad1f9e8),
	.w1(32'hbaaa00e1),
	.w2(32'hba86e721),
	.w3(32'hbabae4e1),
	.w4(32'hba8b37b0),
	.w5(32'h3ac0ecc1),
	.w6(32'hba8da444),
	.w7(32'hbb489d32),
	.w8(32'hb8301d43),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad8c931),
	.w1(32'h38ee3d33),
	.w2(32'hb9319f4b),
	.w3(32'h3a4b0e8b),
	.w4(32'h380bceac),
	.w5(32'h3a77036a),
	.w6(32'hb94e7015),
	.w7(32'h3a259a3e),
	.w8(32'h399dd5eb),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1ada69),
	.w1(32'hb82cfacb),
	.w2(32'h3a3305f1),
	.w3(32'hb9bc5244),
	.w4(32'h3abeed5b),
	.w5(32'h3b734cfa),
	.w6(32'hba245ea3),
	.w7(32'h39ffd3f3),
	.w8(32'h3a6a821e),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2a003a),
	.w1(32'hba2ad25a),
	.w2(32'h3993ed1f),
	.w3(32'h3b67b4f5),
	.w4(32'h3b0c3dce),
	.w5(32'h393880ce),
	.w6(32'h3a013c14),
	.w7(32'h3ac24d12),
	.w8(32'hba5905f4),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98bef96),
	.w1(32'h3a410818),
	.w2(32'h3a6e7e39),
	.w3(32'hb9be324c),
	.w4(32'hb9b6c389),
	.w5(32'h3a543ebf),
	.w6(32'h39ed3438),
	.w7(32'hb996ba37),
	.w8(32'hb90cbcaa),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba96a0bd),
	.w1(32'hba54dc82),
	.w2(32'h39f64329),
	.w3(32'hb9e7dbf5),
	.w4(32'hba589d1b),
	.w5(32'hbab3e335),
	.w6(32'h3923d17f),
	.w7(32'hb950eafe),
	.w8(32'hbb8559c7),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc19e450),
	.w1(32'hbbbbb1b4),
	.w2(32'hba93ce05),
	.w3(32'hbb805dde),
	.w4(32'hbb299e75),
	.w5(32'hb917d50b),
	.w6(32'hbbe4e1c7),
	.w7(32'hbb7db7ab),
	.w8(32'hbaa74940),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaf110a),
	.w1(32'hbb4d2dd7),
	.w2(32'hbb3021b3),
	.w3(32'hbb99449e),
	.w4(32'hbb37905d),
	.w5(32'hba8bb3ad),
	.w6(32'hbb8a7e43),
	.w7(32'hbb52d895),
	.w8(32'hbaea095d),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb90b208),
	.w1(32'hbbb7565b),
	.w2(32'hbbd4ad58),
	.w3(32'hbb995841),
	.w4(32'hbb81539a),
	.w5(32'hbbb3de5f),
	.w6(32'hbb65e18c),
	.w7(32'hbba987d6),
	.w8(32'hbb8649c4),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7b2cd2),
	.w1(32'h3ac28756),
	.w2(32'h3aae6b05),
	.w3(32'h3a899500),
	.w4(32'h3b2f9c73),
	.w5(32'h3aa84268),
	.w6(32'hb98c1b05),
	.w7(32'h391f27ca),
	.w8(32'h3a563414),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8f89dc),
	.w1(32'h3a9f4ee9),
	.w2(32'hbaf66e00),
	.w3(32'h3aa1039c),
	.w4(32'hb9546e97),
	.w5(32'h3a67c722),
	.w6(32'h391d2eac),
	.w7(32'h3b0a0fcb),
	.w8(32'hba2546e3),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8994a9),
	.w1(32'hbbb63a5e),
	.w2(32'hbbbd6417),
	.w3(32'hbaad5fe7),
	.w4(32'hbb4c172d),
	.w5(32'hbb2fdff9),
	.w6(32'hba025edd),
	.w7(32'hbb60ec82),
	.w8(32'hbb0c4e17),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa655e2),
	.w1(32'hbad8ea61),
	.w2(32'hbae8a89c),
	.w3(32'hbb7a6738),
	.w4(32'hbb34f243),
	.w5(32'h3aba5ca3),
	.w6(32'hbb4f2181),
	.w7(32'hba899193),
	.w8(32'h3ae4fe35),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aecf2dd),
	.w1(32'h3b19b813),
	.w2(32'h3a432c11),
	.w3(32'h3a07c883),
	.w4(32'h3a83ca6a),
	.w5(32'hb80cc920),
	.w6(32'h3a49a727),
	.w7(32'h3a99dfb2),
	.w8(32'h3a4eaa2a),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a981aca),
	.w1(32'hbb2c887e),
	.w2(32'hbb7359d1),
	.w3(32'hbafe0904),
	.w4(32'hbb06614d),
	.w5(32'hbabb45a7),
	.w6(32'hba5b7798),
	.w7(32'hbb08eb0a),
	.w8(32'hbae2a7fe),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9972c7e),
	.w1(32'h3a0e5a52),
	.w2(32'h3a246646),
	.w3(32'hb99a2285),
	.w4(32'h3a10f07a),
	.w5(32'hba3e0a51),
	.w6(32'hba194986),
	.w7(32'hba205939),
	.w8(32'hbb180584),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbae0f45),
	.w1(32'hbbb2ab87),
	.w2(32'hbb678f62),
	.w3(32'hbb08dbb5),
	.w4(32'hbb3082a1),
	.w5(32'hba6528c9),
	.w6(32'hbaf89385),
	.w7(32'hbb12f52b),
	.w8(32'h3a73fcbf),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba06d214),
	.w1(32'hbb7fb829),
	.w2(32'hbb53b53d),
	.w3(32'hbadb8dd1),
	.w4(32'hbb01c672),
	.w5(32'hbb793f70),
	.w6(32'hba2d749c),
	.w7(32'hbb1e86b9),
	.w8(32'hbb0bf9d5),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a7c478),
	.w1(32'hb9c07bfd),
	.w2(32'h39f326aa),
	.w3(32'hbadaccd1),
	.w4(32'hb968aa8e),
	.w5(32'h3a7b740a),
	.w6(32'h3ac940b1),
	.w7(32'h3958b065),
	.w8(32'h3ae5b512),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae6cba8),
	.w1(32'hbb3ae235),
	.w2(32'hbacbb403),
	.w3(32'hbae2e6ee),
	.w4(32'hbb33f165),
	.w5(32'h38ca67e1),
	.w6(32'hba6d8c2c),
	.w7(32'hbb1c6900),
	.w8(32'h39c2ca3d),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cd4a4b),
	.w1(32'h3a916e64),
	.w2(32'h3adefbbc),
	.w3(32'hb9da260b),
	.w4(32'h3a5f3376),
	.w5(32'h3b218fbd),
	.w6(32'hba3312c9),
	.w7(32'h3abf2c5f),
	.w8(32'h3b1cda84),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a90c0a3),
	.w1(32'hba92d91c),
	.w2(32'hbaf509e8),
	.w3(32'h3ab037bb),
	.w4(32'hb80dbee9),
	.w5(32'hba05aa16),
	.w6(32'h3b0e24ce),
	.w7(32'h3ac43fef),
	.w8(32'hbab31568),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb28681a),
	.w1(32'hbbb10b3c),
	.w2(32'hbbde986b),
	.w3(32'hbb6a71cc),
	.w4(32'hbaf9a17a),
	.w5(32'hbbd548b5),
	.w6(32'hbb9574eb),
	.w7(32'hbb8252af),
	.w8(32'hbb8c5938),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4a8eee),
	.w1(32'hba1bb902),
	.w2(32'hbb5be6c0),
	.w3(32'hbac15aa2),
	.w4(32'h3a1ddbed),
	.w5(32'hbaa2ee35),
	.w6(32'hbacc760a),
	.w7(32'hbab2499e),
	.w8(32'h3946f080),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b06407f),
	.w1(32'h3af8f3de),
	.w2(32'h3aa1844b),
	.w3(32'h39c3b79e),
	.w4(32'h39bc8187),
	.w5(32'hb9f264c5),
	.w6(32'h3b36c5be),
	.w7(32'h3aadfd7a),
	.w8(32'hba411b55),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba11d981),
	.w1(32'h3a0ee0ee),
	.w2(32'h3a0b31d2),
	.w3(32'h3a966812),
	.w4(32'h3aea1b39),
	.w5(32'h3985ab4c),
	.w6(32'h39d6755d),
	.w7(32'h3a9a8abc),
	.w8(32'hba99b318),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa91548),
	.w1(32'h3953887f),
	.w2(32'hba559e7d),
	.w3(32'hba9866ee),
	.w4(32'hb91c8f50),
	.w5(32'h3b014b84),
	.w6(32'hba6fbe29),
	.w7(32'h38e0d886),
	.w8(32'h3b61e5f0),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b40cf1c),
	.w1(32'h3b0bb210),
	.w2(32'h39a26929),
	.w3(32'h3b03c236),
	.w4(32'h3b6c3c89),
	.w5(32'h3b375e08),
	.w6(32'h3b701b5c),
	.w7(32'h3b8af751),
	.w8(32'h3b287714),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf3d4ab),
	.w1(32'hbb7effdf),
	.w2(32'hbb504bf0),
	.w3(32'hbb8875c8),
	.w4(32'hbb1276ea),
	.w5(32'hbb8e517f),
	.w6(32'hbb52c5c1),
	.w7(32'hbb168ca0),
	.w8(32'hbb300044),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a98b2a1),
	.w1(32'h3a2d528a),
	.w2(32'hb8cd1074),
	.w3(32'hbb14ee0b),
	.w4(32'hbb0b3746),
	.w5(32'h3a375011),
	.w6(32'h3b3ad4be),
	.w7(32'h3a0c37d5),
	.w8(32'hbaba5dae),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb91d313),
	.w1(32'hbb5fbec1),
	.w2(32'hbb2ee687),
	.w3(32'h3b478f5d),
	.w4(32'h3ac9a11b),
	.w5(32'hbb4d96b4),
	.w6(32'h3ae82010),
	.w7(32'h39faeba4),
	.w8(32'h39c66553),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f2603),
	.w1(32'hbb856da0),
	.w2(32'hbaf0bae6),
	.w3(32'hbb43d99e),
	.w4(32'hbb09798f),
	.w5(32'hbb23b8a0),
	.w6(32'hba8d11e1),
	.w7(32'hba182e45),
	.w8(32'hbb7d0a90),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb78e8de),
	.w1(32'hbb635692),
	.w2(32'hbb7424cb),
	.w3(32'hbb483d8b),
	.w4(32'hbb4c2e25),
	.w5(32'hbb107906),
	.w6(32'hbb45d673),
	.w7(32'hbb62ccc1),
	.w8(32'hbaf8d1c9),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa778df),
	.w1(32'hbaa3181c),
	.w2(32'hb93ebfa4),
	.w3(32'hbad071de),
	.w4(32'h39c21442),
	.w5(32'hb6bd9233),
	.w6(32'h39e19bae),
	.w7(32'hba27e590),
	.w8(32'h385860ab),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3085c9),
	.w1(32'hbae53fd5),
	.w2(32'h38073862),
	.w3(32'h38047c1a),
	.w4(32'hbace3550),
	.w5(32'hbb2ef966),
	.w6(32'h390095bd),
	.w7(32'h394e97ce),
	.w8(32'h3b1d313d),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d01702),
	.w1(32'hbafd684c),
	.w2(32'hbb2ac199),
	.w3(32'hbb8d3e95),
	.w4(32'hbbc5c1a7),
	.w5(32'hbb4ef2e7),
	.w6(32'h3b07a53e),
	.w7(32'h38ffe7b3),
	.w8(32'hba07db6e),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b110e7d),
	.w1(32'h3bd68827),
	.w2(32'h3b5b50fc),
	.w3(32'h39eab1b9),
	.w4(32'h3c016e47),
	.w5(32'h3bd1e894),
	.w6(32'hbb1df7c8),
	.w7(32'h3bb5b6e4),
	.w8(32'h3b9c0ab3),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb891fca8),
	.w1(32'h3bc40abe),
	.w2(32'h3bb4b7e6),
	.w3(32'h3b8c0699),
	.w4(32'h3c27f5f9),
	.w5(32'h3b262a47),
	.w6(32'h3b943662),
	.w7(32'h3c18e662),
	.w8(32'h3b84fb15),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaea2d34),
	.w1(32'hba23c8e5),
	.w2(32'hbabefbcc),
	.w3(32'hbb2fdeb3),
	.w4(32'hba94356e),
	.w5(32'hb9828d20),
	.w6(32'hbb8f29cf),
	.w7(32'hbab4ca59),
	.w8(32'h39bb384e),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1644e6),
	.w1(32'hba20dae4),
	.w2(32'hbad638d1),
	.w3(32'hba574fe7),
	.w4(32'hba6ee06a),
	.w5(32'h3a8719ea),
	.w6(32'hbacbef40),
	.w7(32'hbab80520),
	.w8(32'h3ab31649),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f4492c),
	.w1(32'h3a2138ea),
	.w2(32'h3a3ca651),
	.w3(32'h3a8b0627),
	.w4(32'h3a7f8052),
	.w5(32'hba5905bd),
	.w6(32'h3aef92fa),
	.w7(32'h3b0ab838),
	.w8(32'hba87862c),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6ff734),
	.w1(32'hbb3f9c30),
	.w2(32'hbb255fab),
	.w3(32'hb93c4c9f),
	.w4(32'h3b01d868),
	.w5(32'hb9c844fc),
	.w6(32'hb9b48877),
	.w7(32'h3a32760f),
	.w8(32'hbad90c6d),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc01cfbf),
	.w1(32'hbbaeaba8),
	.w2(32'hbbbee4fd),
	.w3(32'hbc01063b),
	.w4(32'hbae2f3d3),
	.w5(32'hbbf63d83),
	.w6(32'hba733e19),
	.w7(32'hba9bbf61),
	.w8(32'hbb838bc8),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc11e5df),
	.w1(32'hbc0cfe06),
	.w2(32'hbc01e9a2),
	.w3(32'hbc15102f),
	.w4(32'hbbf1998d),
	.w5(32'hba087637),
	.w6(32'hbc0664e7),
	.w7(32'hbbb9c83d),
	.w8(32'hba38cdbd),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb43d4de),
	.w1(32'hbb5e2ac9),
	.w2(32'hbbaa0d81),
	.w3(32'hb9df597d),
	.w4(32'hba5a9e0b),
	.w5(32'hbb48401c),
	.w6(32'h3901f054),
	.w7(32'hba6d1e99),
	.w8(32'hbb7a9ec6),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc26715b),
	.w1(32'hbc0f4de8),
	.w2(32'hbbf83e5e),
	.w3(32'hbc0ea61d),
	.w4(32'hbbd0b050),
	.w5(32'hbbb1c342),
	.w6(32'hbbedcc9d),
	.w7(32'hbba68b54),
	.w8(32'hbba6eb19),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb08744e),
	.w1(32'hbb9d431b),
	.w2(32'hbb905d9b),
	.w3(32'hb88f38ec),
	.w4(32'hbb58406b),
	.w5(32'hbbacb951),
	.w6(32'h3a89ae33),
	.w7(32'hbb0e9783),
	.w8(32'hbba086d2),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5270fc),
	.w1(32'hbb45dbc0),
	.w2(32'hbb9340cf),
	.w3(32'hbabaf249),
	.w4(32'hb9d47bf4),
	.w5(32'h3a6faaea),
	.w6(32'hbac6970d),
	.w7(32'hbaecd74b),
	.w8(32'h3a787e29),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b0f645),
	.w1(32'h3a300899),
	.w2(32'h3abe9c8e),
	.w3(32'hb9e7c0f6),
	.w4(32'hba08369d),
	.w5(32'hbab28678),
	.w6(32'hba60c722),
	.w7(32'hb93edb68),
	.w8(32'hbb4ca0a9),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b29fc32),
	.w1(32'h3b197ce7),
	.w2(32'h3a4eef51),
	.w3(32'h3b415d9f),
	.w4(32'h3b02d825),
	.w5(32'h3aa7c16f),
	.w6(32'h3b1d92f3),
	.w7(32'h3b205539),
	.w8(32'h3823a477),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e0799c),
	.w1(32'hb9b7ac2b),
	.w2(32'hba4871df),
	.w3(32'h3ae875db),
	.w4(32'h3b0e8301),
	.w5(32'hba194e1f),
	.w6(32'h3a68cd0d),
	.w7(32'h39a36a2f),
	.w8(32'hba950f05),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ba29a7),
	.w1(32'hb9ee19c9),
	.w2(32'hba50d2ce),
	.w3(32'hba73409b),
	.w4(32'hba970fc9),
	.w5(32'hbab34863),
	.w6(32'hba2aba27),
	.w7(32'hba1f880c),
	.w8(32'h3a6246e2),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad73e32),
	.w1(32'hba9511e3),
	.w2(32'hbb9e3428),
	.w3(32'hba889f4a),
	.w4(32'hbb4e8cb9),
	.w5(32'hbb597c9d),
	.w6(32'h3a81c350),
	.w7(32'hbaaa3e87),
	.w8(32'hbb2f1918),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba32beba),
	.w1(32'hbacd6f10),
	.w2(32'hba87b30c),
	.w3(32'h354802a8),
	.w4(32'h39bcab1d),
	.w5(32'hba576775),
	.w6(32'h3a0640f1),
	.w7(32'hba18bf6d),
	.w8(32'hba33042f),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab71957),
	.w1(32'hbad8ba40),
	.w2(32'hbad0af5e),
	.w3(32'hbad01ce1),
	.w4(32'h39153643),
	.w5(32'hbb0dee55),
	.w6(32'hbafda1a1),
	.w7(32'hbae3dddc),
	.w8(32'h383ecbba),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aae45c8),
	.w1(32'hb9c48d0b),
	.w2(32'hbad905c5),
	.w3(32'hba19391e),
	.w4(32'hb7159691),
	.w5(32'h3a4b403a),
	.w6(32'hb9ef7b30),
	.w7(32'hba3157a3),
	.w8(32'h3a9393f9),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a75ad4e),
	.w1(32'h399c0d28),
	.w2(32'h3a46f22c),
	.w3(32'hb9cf3b60),
	.w4(32'hba0d7b25),
	.w5(32'h3af6d1f4),
	.w6(32'h3a8eca64),
	.w7(32'h381baca2),
	.w8(32'h3a92dc1c),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a37e0cb),
	.w1(32'h3ac63803),
	.w2(32'h3b2c8f09),
	.w3(32'h3abf90df),
	.w4(32'h3b15c3f6),
	.w5(32'h3af09a27),
	.w6(32'hba1a9941),
	.w7(32'h3b0ebc3d),
	.w8(32'h3adae5b6),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a55ab4),
	.w1(32'h3aeff21d),
	.w2(32'h3a7afcee),
	.w3(32'h3af54542),
	.w4(32'h3b120a64),
	.w5(32'h3b980b23),
	.w6(32'h3a6b1703),
	.w7(32'h3aaf3b08),
	.w8(32'h3aef46c0),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0943d9),
	.w1(32'h396a6f01),
	.w2(32'h3ad0deb9),
	.w3(32'h3b1981ff),
	.w4(32'h3b702afe),
	.w5(32'h3ab526ef),
	.w6(32'h3b05ed14),
	.w7(32'h3b73c822),
	.w8(32'h3ae47676),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a01c41f),
	.w1(32'h3ae75bef),
	.w2(32'h3abf8291),
	.w3(32'h3a4d5dd9),
	.w4(32'h3b2a5ed1),
	.w5(32'h39086bec),
	.w6(32'h3b58fd9c),
	.w7(32'h3ad6971b),
	.w8(32'hb8d5fd16),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb074f48),
	.w1(32'hbb0379d4),
	.w2(32'h38274889),
	.w3(32'hba9c9869),
	.w4(32'h3a5ff722),
	.w5(32'h39b7131c),
	.w6(32'hb97a660a),
	.w7(32'h3a052fbd),
	.w8(32'h3a61e277),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1fa85d),
	.w1(32'hb7ae6635),
	.w2(32'hba3795ba),
	.w3(32'hb5239cc4),
	.w4(32'h398afd00),
	.w5(32'hbad1c389),
	.w6(32'hb978dc0a),
	.w7(32'hba665f83),
	.w8(32'hb9b549b0),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac2c455),
	.w1(32'hba3b9063),
	.w2(32'h3ad0f5cc),
	.w3(32'hb9ab1171),
	.w4(32'h3aa11d70),
	.w5(32'h39bafefd),
	.w6(32'h3ab3e84d),
	.w7(32'h3abc85a5),
	.w8(32'hbb1e3e75),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaed7a13),
	.w1(32'hbb1706a5),
	.w2(32'hbac7ad0f),
	.w3(32'hb942ee94),
	.w4(32'hba8239a9),
	.w5(32'h3ab43407),
	.w6(32'hba7550ba),
	.w7(32'hbb176c22),
	.w8(32'h3a901fa3),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac0a050),
	.w1(32'hbacba825),
	.w2(32'hbaf7b0fd),
	.w3(32'hbb3364cb),
	.w4(32'hbb51a487),
	.w5(32'hbb73e62f),
	.w6(32'h3a461a6d),
	.w7(32'h38a0e448),
	.w8(32'hb9ff9029),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb717402),
	.w1(32'hb9a20798),
	.w2(32'hbb0f662a),
	.w3(32'hbb88d50e),
	.w4(32'hbb0e504c),
	.w5(32'hbb1aabbc),
	.w6(32'hbb0c5b34),
	.w7(32'hbb4b794b),
	.w8(32'hbb275b3a),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb340a38),
	.w1(32'h38b6feb5),
	.w2(32'h39ce3d60),
	.w3(32'hbabb2a99),
	.w4(32'h3b1d2fcd),
	.w5(32'h3ada3f3b),
	.w6(32'h39e60b7f),
	.w7(32'h3b032537),
	.w8(32'h3a379526),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb890118),
	.w1(32'hba97fe1a),
	.w2(32'hbbd1a32e),
	.w3(32'hbb8412fa),
	.w4(32'hba923406),
	.w5(32'hbbc6d8af),
	.w6(32'hbb329bb8),
	.w7(32'hbb2995ed),
	.w8(32'hbb955bf7),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb984e7ab),
	.w1(32'hba2030fd),
	.w2(32'hb844f191),
	.w3(32'hb9b0b03c),
	.w4(32'hb85dcd1b),
	.w5(32'h3aeefce2),
	.w6(32'h3a381952),
	.w7(32'hb7d394ca),
	.w8(32'h3a1ab1f0),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d298a8),
	.w1(32'hb95f68e0),
	.w2(32'h3ad9db7c),
	.w3(32'h39929da8),
	.w4(32'hba0fae5b),
	.w5(32'hbaa7ce72),
	.w6(32'hb933563c),
	.w7(32'hb947d99c),
	.w8(32'h3b35b53f),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f51afa),
	.w1(32'h3a831ef1),
	.w2(32'h3a01b2d6),
	.w3(32'hba8b01ac),
	.w4(32'h3a2e37b2),
	.w5(32'hbb3e38e7),
	.w6(32'h3b494b81),
	.w7(32'h3aee889b),
	.w8(32'hbb305bb9),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb47ea2c),
	.w1(32'hbb585251),
	.w2(32'hbb00d6b6),
	.w3(32'hbb180d6e),
	.w4(32'hbae5b4f6),
	.w5(32'hb8a1150e),
	.w6(32'hbabf22ed),
	.w7(32'hba8e96c1),
	.w8(32'h3a46a146),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acd415d),
	.w1(32'h3a8ddf8d),
	.w2(32'h3a1706fe),
	.w3(32'hba42d7f2),
	.w4(32'hbaf78898),
	.w5(32'hbb252543),
	.w6(32'h3a8315ab),
	.w7(32'hbab1a11b),
	.w8(32'hbb475549),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5575df),
	.w1(32'hbb5536fe),
	.w2(32'hbb372ea7),
	.w3(32'hbb3256b3),
	.w4(32'hbb4da2f9),
	.w5(32'h3b121317),
	.w6(32'hbb11d7eb),
	.w7(32'hbb2541b8),
	.w8(32'h3ae9ae1b),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf25950),
	.w1(32'hbae38875),
	.w2(32'hbabdaf57),
	.w3(32'hba3d7fd2),
	.w4(32'hbaa11716),
	.w5(32'hba05b397),
	.w6(32'hbb1dcb9c),
	.w7(32'hba29fbf4),
	.w8(32'hbaeb8f54),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9acde1e),
	.w1(32'hbb8fea5f),
	.w2(32'hbba91d9d),
	.w3(32'hbacf2c65),
	.w4(32'hbb8899e5),
	.w5(32'hbb553943),
	.w6(32'hbb43bb12),
	.w7(32'hbb608471),
	.w8(32'hbb3a4bef),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba98d27a),
	.w1(32'h3a8f897b),
	.w2(32'h36c28f13),
	.w3(32'h39faf3ae),
	.w4(32'h39086edf),
	.w5(32'h39fedca2),
	.w6(32'hb95ef873),
	.w7(32'h3a8ca91e),
	.w8(32'hba8a549c),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ad6a57),
	.w1(32'hb90afd7d),
	.w2(32'hba9224b1),
	.w3(32'hb9fb2960),
	.w4(32'hbab6ab24),
	.w5(32'hbb9c523f),
	.w6(32'h3a601bac),
	.w7(32'hbabbdc33),
	.w8(32'hbbac3924),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd46c51),
	.w1(32'hbba745bf),
	.w2(32'hbb8f4386),
	.w3(32'hbba23db5),
	.w4(32'hbb8fe3f6),
	.w5(32'hbb787eb0),
	.w6(32'hbbf233f9),
	.w7(32'hbb85e6ba),
	.w8(32'hbb7f08ef),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb471954),
	.w1(32'hbba10e0c),
	.w2(32'hbba1d8c6),
	.w3(32'hbb25c899),
	.w4(32'hbb68b61f),
	.w5(32'hb815f29d),
	.w6(32'hbb004cd5),
	.w7(32'hbb1b781e),
	.w8(32'hb93c1b3a),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb850a7da),
	.w1(32'h3906ebdc),
	.w2(32'h39d4bf0d),
	.w3(32'h3a8076b0),
	.w4(32'h39f292d0),
	.w5(32'hba6adde2),
	.w6(32'hb9c28b4f),
	.w7(32'h3a1f859d),
	.w8(32'h3b07a49b),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1ef42b),
	.w1(32'h3ae60496),
	.w2(32'h39e53692),
	.w3(32'hb930621f),
	.w4(32'hb6991416),
	.w5(32'h3a21c1c6),
	.w6(32'h3aac65b2),
	.w7(32'h39dc5cd0),
	.w8(32'hb84c7f2d),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb92d6033),
	.w1(32'hba3a6fcc),
	.w2(32'hb9483b8c),
	.w3(32'h39b4f07f),
	.w4(32'hba898ff5),
	.w5(32'h3b8154a7),
	.w6(32'hba851aed),
	.w7(32'hba4c8205),
	.w8(32'h3ad6d669),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d1f6d4),
	.w1(32'h3a3e1ff5),
	.w2(32'h3a28f189),
	.w3(32'h3b09a310),
	.w4(32'h3ae626c1),
	.w5(32'h39c510a1),
	.w6(32'h3b301bed),
	.w7(32'h3a759317),
	.w8(32'h3a2c2324),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1ceea2),
	.w1(32'h3a30c327),
	.w2(32'hbac18176),
	.w3(32'hbaf139fa),
	.w4(32'hba4cb82a),
	.w5(32'hb7ca9eb1),
	.w6(32'hbabd3167),
	.w7(32'hb8559ba0),
	.w8(32'hba9d4bdb),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399cd12b),
	.w1(32'hba3c42df),
	.w2(32'hb8fbd56c),
	.w3(32'hb6ac4a53),
	.w4(32'hba01e231),
	.w5(32'h39a44174),
	.w6(32'hba53fc4c),
	.w7(32'hba943251),
	.w8(32'hba7f7994),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391252d9),
	.w1(32'hb9b327f3),
	.w2(32'hba8a12b8),
	.w3(32'h3a95d73c),
	.w4(32'h39b45ad6),
	.w5(32'hbb1131ff),
	.w6(32'hb9b0ac4e),
	.w7(32'hbabb3ccb),
	.w8(32'hbacd455f),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8b4757),
	.w1(32'h3a5ad18e),
	.w2(32'h3a50b170),
	.w3(32'h3a9ecae5),
	.w4(32'h3ace17ae),
	.w5(32'h3a6fe762),
	.w6(32'h398bd53e),
	.w7(32'h3b0ff358),
	.w8(32'hb9f8fc87),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa25daf),
	.w1(32'hb7cc231a),
	.w2(32'hbb3420df),
	.w3(32'hbad5c629),
	.w4(32'h3ad2c26a),
	.w5(32'h3a6ac52f),
	.w6(32'hbae8ca9a),
	.w7(32'hba05db57),
	.w8(32'h3aa59b78),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb338ee2),
	.w1(32'h3a9b7276),
	.w2(32'hba23c46c),
	.w3(32'hbb2a472e),
	.w4(32'hbb5d1321),
	.w5(32'hbb72adca),
	.w6(32'hb99a4ede),
	.w7(32'h38ee1e64),
	.w8(32'hbb076998),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394055da),
	.w1(32'h39e4c525),
	.w2(32'hb9b2298c),
	.w3(32'h3b19878e),
	.w4(32'h3b06d6a8),
	.w5(32'h3a742d9f),
	.w6(32'h3ae17f03),
	.w7(32'h3ace31fd),
	.w8(32'h39d6c9dc),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb323bea),
	.w1(32'hba1dee97),
	.w2(32'hbb33332f),
	.w3(32'hb99c99d5),
	.w4(32'h39f8d0f8),
	.w5(32'hbab3ce7e),
	.w6(32'hba5e03df),
	.w7(32'hb9a349c2),
	.w8(32'hba15fae6),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab20ebf),
	.w1(32'h39719799),
	.w2(32'h38498dfa),
	.w3(32'h3a10d3b5),
	.w4(32'h38f450ce),
	.w5(32'h3abcf5aa),
	.w6(32'h3abe04db),
	.w7(32'h3ab13fda),
	.w8(32'h3a1936ec),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba27de4a),
	.w1(32'hb9577cec),
	.w2(32'hba956a54),
	.w3(32'h3ab49c7e),
	.w4(32'h3afb0751),
	.w5(32'hbb26a63e),
	.w6(32'hba5c1e18),
	.w7(32'h3a1acd3f),
	.w8(32'hbb33d552),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb317062),
	.w1(32'hb9a70851),
	.w2(32'h3b26fb5b),
	.w3(32'hb98489a7),
	.w4(32'h39e89686),
	.w5(32'hba8efab6),
	.w6(32'h3afcf0d9),
	.w7(32'h3b8ce94a),
	.w8(32'hba0b8484),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8314bd),
	.w1(32'hbb03ec8f),
	.w2(32'hbaf3ee00),
	.w3(32'hbaada68a),
	.w4(32'hb8d8f4cb),
	.w5(32'h3aa9e25c),
	.w6(32'h3a5df910),
	.w7(32'hb9be3c0f),
	.w8(32'h3b24e50b),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b032b71),
	.w1(32'h3c1d6763),
	.w2(32'h3b80ac78),
	.w3(32'h3b84c5bb),
	.w4(32'h39b6e9c7),
	.w5(32'hbb07db45),
	.w6(32'h3bc70119),
	.w7(32'h3b105a69),
	.w8(32'hbbcc4dd3),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1ee567),
	.w1(32'hbb8e83a9),
	.w2(32'hbbf82fa9),
	.w3(32'hbc12f363),
	.w4(32'h39aa4179),
	.w5(32'h3b39141d),
	.w6(32'hbb06b317),
	.w7(32'hbbec0e95),
	.w8(32'h3bb25f39),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc49cba2),
	.w1(32'hbc058644),
	.w2(32'hbc0b9c5b),
	.w3(32'hbc1b994b),
	.w4(32'hbb6024d9),
	.w5(32'h3aa4f578),
	.w6(32'hbc103501),
	.w7(32'hba13997e),
	.w8(32'hbb6ad4e1),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc02021b),
	.w1(32'hbbc102cb),
	.w2(32'hbc3d1c38),
	.w3(32'h3b4c4938),
	.w4(32'hba4cd085),
	.w5(32'hbb8a122c),
	.w6(32'h3a0600f9),
	.w7(32'hbabe3a47),
	.w8(32'hbbb1ead2),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0b1ee9),
	.w1(32'hbaaf5865),
	.w2(32'hb9b81e8c),
	.w3(32'hbc113638),
	.w4(32'hbacd6b6f),
	.w5(32'hbbb9a74e),
	.w6(32'hbbd3a69a),
	.w7(32'h3bbdcd26),
	.w8(32'h3a34fefc),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbef6461),
	.w1(32'hbb05cb4d),
	.w2(32'hbaab7b19),
	.w3(32'hbb9d8ba2),
	.w4(32'h3bade247),
	.w5(32'h3c0898db),
	.w6(32'h3a9d917f),
	.w7(32'h3b63958e),
	.w8(32'h3be8c785),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c7149),
	.w1(32'hba8ff0d6),
	.w2(32'hbc46b61a),
	.w3(32'hbb9a10e5),
	.w4(32'hbba15b4d),
	.w5(32'hbb1fd41a),
	.w6(32'h3acb0927),
	.w7(32'hbc3f8403),
	.w8(32'hbc146999),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5e8934),
	.w1(32'hbb80be4a),
	.w2(32'hbaef7ff0),
	.w3(32'hbbdce282),
	.w4(32'hbb4e9620),
	.w5(32'h3bb547d4),
	.w6(32'hbc1119e2),
	.w7(32'h3b020e04),
	.w8(32'hbb39fd3e),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad334f6),
	.w1(32'hba084d5e),
	.w2(32'hbbc4942d),
	.w3(32'hbaf705b1),
	.w4(32'h3aa9191f),
	.w5(32'hbc68d822),
	.w6(32'hbb27776d),
	.w7(32'h391fe2ad),
	.w8(32'hbb80e711),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbeab649),
	.w1(32'hbb13a077),
	.w2(32'hba6f9f32),
	.w3(32'hbbce288d),
	.w4(32'hbbc11bfc),
	.w5(32'h3a794fb4),
	.w6(32'h3be376c1),
	.w7(32'hbaa431af),
	.w8(32'h3bb73ac7),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abfff3c),
	.w1(32'h3bdb6cd6),
	.w2(32'hbb4eee03),
	.w3(32'h3c3aa9ae),
	.w4(32'hbb313be4),
	.w5(32'hbc766928),
	.w6(32'h3c82a75a),
	.w7(32'h387ddcb9),
	.w8(32'hbc2e8250),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1f3a37),
	.w1(32'h3c1f6769),
	.w2(32'h3c75c126),
	.w3(32'h39133db0),
	.w4(32'h3b8dd0d3),
	.w5(32'hbb5c5e9d),
	.w6(32'h3c43422c),
	.w7(32'h3c3090e5),
	.w8(32'hbc162b80),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1704fa),
	.w1(32'h3b93378a),
	.w2(32'hbb6aa2f9),
	.w3(32'hbab5e9d3),
	.w4(32'h3b4dde81),
	.w5(32'hbaa48b5b),
	.w6(32'h3b2d14b9),
	.w7(32'h3b1d6230),
	.w8(32'hbbba41b5),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc161a55),
	.w1(32'h3ad352e3),
	.w2(32'hbb3c1c41),
	.w3(32'hbb89ccae),
	.w4(32'hbaadce2d),
	.w5(32'h38a03606),
	.w6(32'hbb1555a7),
	.w7(32'hbb34cc8a),
	.w8(32'hbc0e123c),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b43ff08),
	.w1(32'h3c702774),
	.w2(32'h3bbb61fa),
	.w3(32'h3bd1afae),
	.w4(32'h3b9e05f6),
	.w5(32'h3b9154c6),
	.w6(32'h3b59626e),
	.w7(32'h3b35c3df),
	.w8(32'h3b825e42),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb945b4d),
	.w1(32'hbbae817e),
	.w2(32'hbb108f9d),
	.w3(32'hba95f00e),
	.w4(32'hbb7f3515),
	.w5(32'hb9991c83),
	.w6(32'h3b4dff0b),
	.w7(32'h3a9baf9d),
	.w8(32'hbc0856f1),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8bc047),
	.w1(32'h3aee66c6),
	.w2(32'hba85c258),
	.w3(32'h3a62d818),
	.w4(32'hbb8407f0),
	.w5(32'h3b04c33b),
	.w6(32'hbaa035c2),
	.w7(32'hbc08c4a1),
	.w8(32'hbc10eab0),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbed096e),
	.w1(32'h3a578ac9),
	.w2(32'hb97c25fb),
	.w3(32'h3a8fb623),
	.w4(32'hbac64979),
	.w5(32'h3c54d6d9),
	.w6(32'hbb7b14ee),
	.w7(32'hb8344e94),
	.w8(32'h3c0be3d9),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b40ca42),
	.w1(32'hb9505385),
	.w2(32'h3bc3cf97),
	.w3(32'h3c0d3019),
	.w4(32'h3b606c2d),
	.w5(32'hba70c7c9),
	.w6(32'h3b8c1359),
	.w7(32'h3bba59ab),
	.w8(32'h3be0e217),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9fb66f),
	.w1(32'hbb3ec092),
	.w2(32'hbb075215),
	.w3(32'hbba08f97),
	.w4(32'hba3a57bd),
	.w5(32'hbae08d5f),
	.w6(32'hbb1b3943),
	.w7(32'hbbce5c7d),
	.w8(32'h3a9f7dbe),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba553ab),
	.w1(32'hbaa21c13),
	.w2(32'h3a835449),
	.w3(32'hba249e89),
	.w4(32'hbb2e6bf5),
	.w5(32'h3a3e65aa),
	.w6(32'h3ad148a0),
	.w7(32'hb932fab4),
	.w8(32'h3b86cf10),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb982bf7),
	.w1(32'hbaf0f1a2),
	.w2(32'hbbb7944c),
	.w3(32'h3bb6dd7e),
	.w4(32'hb8e0fdf7),
	.w5(32'h3c9defa8),
	.w6(32'h3bb12075),
	.w7(32'h3ada4505),
	.w8(32'h3c103c7b),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3b5a06),
	.w1(32'hbb5df8f8),
	.w2(32'hba0c6796),
	.w3(32'hb98273f7),
	.w4(32'h3b56b359),
	.w5(32'h3c0fdf23),
	.w6(32'hbc2c96c0),
	.w7(32'h3b03dd2c),
	.w8(32'h3bfba253),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf9ce1a),
	.w1(32'h39acfcc9),
	.w2(32'h3c0d0b43),
	.w3(32'hbb828104),
	.w4(32'hbb15dc38),
	.w5(32'h3b4e0be0),
	.w6(32'hbc8e10c4),
	.w7(32'h3c18c76f),
	.w8(32'h3a2d17d2),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c045a6c),
	.w1(32'h3c072f38),
	.w2(32'h3b6c1387),
	.w3(32'h3b963ea6),
	.w4(32'h3c5bfb44),
	.w5(32'h3bd6cb7e),
	.w6(32'hbb8b0345),
	.w7(32'h3bd80f0c),
	.w8(32'hbb9b591a),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2b5cd0),
	.w1(32'h3bcfdc55),
	.w2(32'h3b890dee),
	.w3(32'hba833cf6),
	.w4(32'hbba9eace),
	.w5(32'h391466c4),
	.w6(32'h3926ddc4),
	.w7(32'hb9c789b7),
	.w8(32'h3b3d58e0),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0ca595),
	.w1(32'h3c015049),
	.w2(32'h3ad606f9),
	.w3(32'h3b8af7da),
	.w4(32'hb9c3596e),
	.w5(32'hbb8e01f0),
	.w6(32'h3bb9699c),
	.w7(32'h3c66a500),
	.w8(32'h3be76801),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbda659),
	.w1(32'h3ab7a708),
	.w2(32'h3aa89e07),
	.w3(32'h3ae17f62),
	.w4(32'h3b732e84),
	.w5(32'hbb4c2775),
	.w6(32'h3b1c8e58),
	.w7(32'h3ac8cfcb),
	.w8(32'h3b0d7d22),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8aa61d2),
	.w1(32'h3b9d4821),
	.w2(32'h3bda4ba6),
	.w3(32'h3c191548),
	.w4(32'hbada6f68),
	.w5(32'hbba8040f),
	.w6(32'h3bf781b4),
	.w7(32'h3ba6ce54),
	.w8(32'hbbbbcde4),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9a93e3),
	.w1(32'hbc1ad87e),
	.w2(32'hbb3d994c),
	.w3(32'hb89905b0),
	.w4(32'hbb4068e7),
	.w5(32'hbc025988),
	.w6(32'h3abceb1d),
	.w7(32'hbba8e1d8),
	.w8(32'hbc48e7ab),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b920eff),
	.w1(32'h3c36953e),
	.w2(32'h3c4ddd87),
	.w3(32'hbbb4b5d8),
	.w4(32'h3c240f8b),
	.w5(32'h3b72108f),
	.w6(32'hbacca9e9),
	.w7(32'h3c8b949b),
	.w8(32'hbb0f3ae1),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3232f0),
	.w1(32'hb92f037c),
	.w2(32'h3b05c5ee),
	.w3(32'h3b7259aa),
	.w4(32'hbbc1e699),
	.w5(32'h3bceeaa5),
	.w6(32'hbc262f90),
	.w7(32'hbb6d2c41),
	.w8(32'h3b8f779a),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba51f0a),
	.w1(32'hbbe8f88b),
	.w2(32'hba38c4d4),
	.w3(32'hbaa622d4),
	.w4(32'hbc1e53da),
	.w5(32'h3afb8f2f),
	.w6(32'hbb90e84d),
	.w7(32'hbaf79cb5),
	.w8(32'h3a7df21d),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3939daac),
	.w1(32'hb9a3d1a7),
	.w2(32'hbb65d5aa),
	.w3(32'h3b908ff7),
	.w4(32'hba81a955),
	.w5(32'hbb26ffc7),
	.w6(32'h3b07572a),
	.w7(32'hbb2d623c),
	.w8(32'h3b4e8137),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6c36ef),
	.w1(32'hbba35d5f),
	.w2(32'hbc4c456b),
	.w3(32'hba2800e0),
	.w4(32'hbbbdd7e9),
	.w5(32'hbbca1dc7),
	.w6(32'hba114483),
	.w7(32'hbc1eabe7),
	.w8(32'hbba2d175),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3c7054),
	.w1(32'h3bb4a693),
	.w2(32'h3c0300eb),
	.w3(32'h3a1c2e55),
	.w4(32'h3a88d9b3),
	.w5(32'hb9ec091d),
	.w6(32'h3b81b88d),
	.w7(32'h3c0849f6),
	.w8(32'hbb72b102),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc419e3),
	.w1(32'hba6aaf6c),
	.w2(32'hbb39038a),
	.w3(32'hba61202d),
	.w4(32'hbbc298c0),
	.w5(32'hbbcce4dd),
	.w6(32'hbb21e1ff),
	.w7(32'hb9a1917c),
	.w8(32'h39307ecb),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d72de2),
	.w1(32'hba4b8099),
	.w2(32'hbb60f7d6),
	.w3(32'hba9ec5be),
	.w4(32'h3c014774),
	.w5(32'hba184c78),
	.w6(32'hbba0e513),
	.w7(32'h3affcd4d),
	.w8(32'hbbd56174),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab99771),
	.w1(32'h3be15a90),
	.w2(32'h3c13decf),
	.w3(32'h3af75f1e),
	.w4(32'h3b82659c),
	.w5(32'hbbeb5431),
	.w6(32'h3b1cab35),
	.w7(32'h3c3d5863),
	.w8(32'hbbacc0e8),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb995f10),
	.w1(32'h3b4cc9c6),
	.w2(32'h3c221515),
	.w3(32'hba9030a4),
	.w4(32'hba006908),
	.w5(32'h39732bcf),
	.w6(32'h3b981de5),
	.w7(32'h3c047d7b),
	.w8(32'hbb739120),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc145ab9),
	.w1(32'hbb8c3391),
	.w2(32'hbb9429b0),
	.w3(32'hba5aae98),
	.w4(32'hbb94d2da),
	.w5(32'hbb35d1ad),
	.w6(32'hbbad28d2),
	.w7(32'h3b0db044),
	.w8(32'h3b42964a),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcbc22a),
	.w1(32'hbc16c020),
	.w2(32'hbb2fba64),
	.w3(32'h396bd113),
	.w4(32'hbc0691fe),
	.w5(32'hbc6feb8c),
	.w6(32'hbb8c1a2f),
	.w7(32'h3b15e30a),
	.w8(32'hbc39d12e),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1d90cf),
	.w1(32'hb7e6ca9e),
	.w2(32'h3b348759),
	.w3(32'hbc2849c4),
	.w4(32'h3bf1a16f),
	.w5(32'hbb822330),
	.w6(32'hbbbbd006),
	.w7(32'hbb81923e),
	.w8(32'hbbbc00b2),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a88b822),
	.w1(32'h3aca6a4e),
	.w2(32'hbb9fe844),
	.w3(32'h3a368233),
	.w4(32'hbb786a36),
	.w5(32'hbb89ebc4),
	.w6(32'hbaf11de7),
	.w7(32'hbba2e106),
	.w8(32'hbc04f3e0),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8735f7),
	.w1(32'h3abc0862),
	.w2(32'hbbed173d),
	.w3(32'hbb0466bb),
	.w4(32'hbb5342ad),
	.w5(32'hbc364d7b),
	.w6(32'hbb074ab8),
	.w7(32'hbb3cb2f5),
	.w8(32'hbc0bbcf0),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0bf29a),
	.w1(32'h3b65898d),
	.w2(32'h3954faa0),
	.w3(32'hbb15792c),
	.w4(32'h3ac8d3d7),
	.w5(32'hbc003e81),
	.w6(32'hbbfd447e),
	.w7(32'h3bd9be47),
	.w8(32'hbb6a774a),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba84840),
	.w1(32'h3b00dc29),
	.w2(32'h3b6faa7e),
	.w3(32'hb96e0057),
	.w4(32'hb91166a9),
	.w5(32'h3ac8533b),
	.w6(32'h3b9bc575),
	.w7(32'h39912471),
	.w8(32'hbb181611),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h370d8b97),
	.w1(32'hba9a640e),
	.w2(32'hbb5c5b5d),
	.w3(32'hbb930c5f),
	.w4(32'hbb89dc4c),
	.w5(32'hbb1b1470),
	.w6(32'hbb57e5df),
	.w7(32'hba65c2d9),
	.w8(32'hbac8a113),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38eaffbe),
	.w1(32'h3a6c687f),
	.w2(32'hbbcb376f),
	.w3(32'h39accb3a),
	.w4(32'h3b340926),
	.w5(32'hbb30dca4),
	.w6(32'h39ae137c),
	.w7(32'hb77b1d56),
	.w8(32'h3bbf6867),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b36cf40),
	.w1(32'hbb6b7aec),
	.w2(32'hbc1eae9c),
	.w3(32'hbb9436cc),
	.w4(32'hbb4daf3d),
	.w5(32'hbc25b57b),
	.w6(32'hbb663fde),
	.w7(32'hbb4f6a60),
	.w8(32'hbba4124a),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b178c8f),
	.w1(32'h3b37cc7e),
	.w2(32'h3c622764),
	.w3(32'hbc17cd7f),
	.w4(32'h3c115995),
	.w5(32'h3c1a0903),
	.w6(32'hbc2c9432),
	.w7(32'h3caba0f0),
	.w8(32'h3c109184),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a20ab49),
	.w1(32'hbb42e4fc),
	.w2(32'hbae62c36),
	.w3(32'h3b9fe551),
	.w4(32'hbb371a6d),
	.w5(32'h3b432735),
	.w6(32'h3b5b0f62),
	.w7(32'hbb89728c),
	.w8(32'h39cd6430),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3924cc),
	.w1(32'h3a212252),
	.w2(32'hbb29869d),
	.w3(32'h3a85ff3a),
	.w4(32'hbb23e931),
	.w5(32'hbc8413d3),
	.w6(32'h3a095006),
	.w7(32'h3bab9644),
	.w8(32'hbc6835f5),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba554c10),
	.w1(32'h39c93ba3),
	.w2(32'hba64410e),
	.w3(32'hbbe2c73c),
	.w4(32'hbb1bba42),
	.w5(32'h3a3a3d42),
	.w6(32'h3af06b67),
	.w7(32'h3c16041b),
	.w8(32'hbb826a5a),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad02a0f),
	.w1(32'hbb116cae),
	.w2(32'hbb4c90f7),
	.w3(32'h3c2ab8a8),
	.w4(32'h3b5a7580),
	.w5(32'hbc48699b),
	.w6(32'h3b2d3360),
	.w7(32'h3ac792cc),
	.w8(32'hbb97948e),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf85214),
	.w1(32'h3b718acf),
	.w2(32'hbbdf32d1),
	.w3(32'hbb84124e),
	.w4(32'hbb7b7af1),
	.w5(32'h3bac71ad),
	.w6(32'h3bde22f3),
	.w7(32'hbaaa27fa),
	.w8(32'h3bf10c7e),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af5dd49),
	.w1(32'h3b4743ee),
	.w2(32'hbb1f4131),
	.w3(32'h3c3739c3),
	.w4(32'hb9cea2f0),
	.w5(32'hbb95d6a4),
	.w6(32'h3bffcab1),
	.w7(32'h3932648d),
	.w8(32'hbbe777e4),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbd90c3),
	.w1(32'h3c0586b7),
	.w2(32'h3c64b57e),
	.w3(32'hbbc853ee),
	.w4(32'h3b62cc6c),
	.w5(32'hbc0bd5e1),
	.w6(32'h3a931b5f),
	.w7(32'h3c58580e),
	.w8(32'h399a1ddb),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae97a82),
	.w1(32'h3bbcf0b0),
	.w2(32'h3b9bafe1),
	.w3(32'hba3dc58e),
	.w4(32'h3a5dee8d),
	.w5(32'h3c3f8fed),
	.w6(32'h39fb9fa2),
	.w7(32'h3beb8765),
	.w8(32'h3c089b00),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c215af7),
	.w1(32'h3c301ae4),
	.w2(32'h3bab9633),
	.w3(32'h3a00aacf),
	.w4(32'h3a1fa31a),
	.w5(32'hbb1a4882),
	.w6(32'hbbecd667),
	.w7(32'h3a9642fd),
	.w8(32'hbbefb9f2),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfc80d2),
	.w1(32'hba563d1d),
	.w2(32'h3b311d3f),
	.w3(32'h3ab817d5),
	.w4(32'hbba0266f),
	.w5(32'h3c09f4d6),
	.w6(32'h3ae20e0d),
	.w7(32'hbb172f31),
	.w8(32'hbbaa8df3),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb03897),
	.w1(32'hbb1eb7e0),
	.w2(32'h3ba39c04),
	.w3(32'h3b8caada),
	.w4(32'h3a0e2b83),
	.w5(32'hbbb95d00),
	.w6(32'h3babfaef),
	.w7(32'h3accb4a9),
	.w8(32'hbbde6123),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe04d18),
	.w1(32'hbc194bd5),
	.w2(32'hbc2ad330),
	.w3(32'hbba30ac0),
	.w4(32'h39f7d0dd),
	.w5(32'hbbc238ed),
	.w6(32'hbc076cae),
	.w7(32'hbc04411b),
	.w8(32'hbbe2e9c6),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3b6903),
	.w1(32'hbc079a2f),
	.w2(32'hb9e70e33),
	.w3(32'hbc357f10),
	.w4(32'hbb724151),
	.w5(32'h3b2944a6),
	.w6(32'hbbf58ac9),
	.w7(32'hb85f831b),
	.w8(32'h3b817478),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aeb67f5),
	.w1(32'hbb3d7008),
	.w2(32'hba11f0a6),
	.w3(32'hba96c9b9),
	.w4(32'h3b3fc46a),
	.w5(32'h3a5e651f),
	.w6(32'hbaa09c75),
	.w7(32'h3a9b75fd),
	.w8(32'hbbb719e7),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e3d6fa),
	.w1(32'hbb1ff7ab),
	.w2(32'hbb8ca0c3),
	.w3(32'hbb9e3fc4),
	.w4(32'h3b204164),
	.w5(32'h3a001c34),
	.w6(32'hbc2fd41d),
	.w7(32'h3baa1cc2),
	.w8(32'h3c330437),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b924b94),
	.w1(32'h396fe281),
	.w2(32'hbb91bf0d),
	.w3(32'hb94d6ee3),
	.w4(32'h3aedcf9f),
	.w5(32'h3b725065),
	.w6(32'h3aa6a718),
	.w7(32'hbb6cfb8a),
	.w8(32'hbb773408),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb7d06c),
	.w1(32'h3b51021e),
	.w2(32'hbbe049e4),
	.w3(32'h3ac0e80c),
	.w4(32'hbb9cfbcb),
	.w5(32'h3c30b543),
	.w6(32'hbc11ef73),
	.w7(32'hbb9cd4d7),
	.w8(32'h3b98d078),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h395d9d6d),
	.w1(32'h3b8a153a),
	.w2(32'hbb1f91a1),
	.w3(32'h3bdf211d),
	.w4(32'h3ba98182),
	.w5(32'hbb8b7728),
	.w6(32'h3bd7f20e),
	.w7(32'h3c278a2c),
	.w8(32'hbaa810d7),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5d68ec),
	.w1(32'hbbe9520b),
	.w2(32'hbc5ab478),
	.w3(32'hbbc8d949),
	.w4(32'hbbd51e32),
	.w5(32'hbac86f4d),
	.w6(32'h3a737ead),
	.w7(32'hbc48a515),
	.w8(32'hbb06e0bb),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe78048),
	.w1(32'hbc27556c),
	.w2(32'hbb91b192),
	.w3(32'hbba43e46),
	.w4(32'hbbb7106e),
	.w5(32'hbc3e6d56),
	.w6(32'hbc395cda),
	.w7(32'hbb0d399e),
	.w8(32'hbaca8d21),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9aee04),
	.w1(32'hbb669ac4),
	.w2(32'hbc02c553),
	.w3(32'hbac435e3),
	.w4(32'hbc14d9b9),
	.w5(32'h3c32981a),
	.w6(32'h3b31e61f),
	.w7(32'hbb13a2aa),
	.w8(32'hb94b6d0f),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3afd38a7),
	.w1(32'hba006017),
	.w2(32'hbba7a5ca),
	.w3(32'h3b689ab9),
	.w4(32'h3b266d3b),
	.w5(32'h3b9c4af7),
	.w6(32'hbbd75297),
	.w7(32'h3bfac61e),
	.w8(32'hbb2d559d),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a768f66),
	.w1(32'hbc1c2759),
	.w2(32'hbc03bbbd),
	.w3(32'hbb590608),
	.w4(32'hbc4ab886),
	.w5(32'h3b2044fa),
	.w6(32'hbbcaaf72),
	.w7(32'hbbd1ba9f),
	.w8(32'h3bc3f124),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5b36c6),
	.w1(32'hbc39b0cb),
	.w2(32'hbc2dcff7),
	.w3(32'hbb4bf060),
	.w4(32'hbb911dd8),
	.w5(32'hbc7f1fe7),
	.w6(32'hbaa67322),
	.w7(32'hbbb4af22),
	.w8(32'hb970545a),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5af542),
	.w1(32'hbb3fde39),
	.w2(32'h3c436f70),
	.w3(32'h396de68d),
	.w4(32'hbb3f4179),
	.w5(32'hbb93c024),
	.w6(32'h3c7e41f5),
	.w7(32'h3be83783),
	.w8(32'h3830fa05),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0520f1),
	.w1(32'hbc109240),
	.w2(32'hbc03fddc),
	.w3(32'hbc0704d8),
	.w4(32'hbbbef8f8),
	.w5(32'h3b9bd37a),
	.w6(32'hbbd60c31),
	.w7(32'hbbe599fa),
	.w8(32'h3afd7da7),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba77c51),
	.w1(32'h3c56ede0),
	.w2(32'h3c564b55),
	.w3(32'h3c31af7f),
	.w4(32'h3c3dd06f),
	.w5(32'hbbbb0718),
	.w6(32'h3c0c653f),
	.w7(32'h3c4e2802),
	.w8(32'hbc02c423),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbc2de8),
	.w1(32'hbb88b52d),
	.w2(32'hbbf9e92a),
	.w3(32'hbc4f31d3),
	.w4(32'hbaf30378),
	.w5(32'h3bc6e3f8),
	.w6(32'hbbd6f40c),
	.w7(32'hbaba8d7f),
	.w8(32'h3bb3e8ec),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af76b5b),
	.w1(32'h3bd79e06),
	.w2(32'hbaeb01ae),
	.w3(32'h3c1bbfde),
	.w4(32'hbb45f6df),
	.w5(32'h3c00a5de),
	.w6(32'h3bc8dd97),
	.w7(32'hbb2de8c0),
	.w8(32'h3bf05466),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb37141),
	.w1(32'hbb16412a),
	.w2(32'h3a4092e1),
	.w3(32'hb9c5b865),
	.w4(32'h3b71fd85),
	.w5(32'h3a51d27c),
	.w6(32'hbbbaafe7),
	.w7(32'h3b1ee6e0),
	.w8(32'h3b7de301),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abb4260),
	.w1(32'h3b345a63),
	.w2(32'h3b89cabe),
	.w3(32'h392f8c3e),
	.w4(32'hb9c581f7),
	.w5(32'h3c004e54),
	.w6(32'h3b9bb3bd),
	.w7(32'h3bc1448c),
	.w8(32'h3b4c77a3),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc22c639),
	.w1(32'hbc2c8ed5),
	.w2(32'hbc0058bb),
	.w3(32'hbb2a1644),
	.w4(32'h3b196663),
	.w5(32'h3c1ee99c),
	.w6(32'hbbf56c39),
	.w7(32'h3b2a06f8),
	.w8(32'h3c99b2d3),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c356845),
	.w1(32'h3b707487),
	.w2(32'h3bf71742),
	.w3(32'hbbaaaa0f),
	.w4(32'hbba546c1),
	.w5(32'hbac32c56),
	.w6(32'hbbe624d8),
	.w7(32'h3b711f9f),
	.w8(32'h3b80208e),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac87f93),
	.w1(32'h3b21e4a7),
	.w2(32'hba65c822),
	.w3(32'h3adf3816),
	.w4(32'hbb03bfc6),
	.w5(32'hbb0e8366),
	.w6(32'h3b86f012),
	.w7(32'h39f63f2b),
	.w8(32'hbaa5a7d2),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9bd320),
	.w1(32'h3b47dbaf),
	.w2(32'h3bf10ccc),
	.w3(32'h3b014c84),
	.w4(32'hbb4f554e),
	.w5(32'hbaa829d0),
	.w6(32'hb9a20979),
	.w7(32'h3b4f6f2a),
	.w8(32'hbb9a6c65),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a70f7a7),
	.w1(32'hbada0e9e),
	.w2(32'h399c534c),
	.w3(32'h3b8c774e),
	.w4(32'h3a9f37f7),
	.w5(32'h3b20860a),
	.w6(32'h3b5467a3),
	.w7(32'hb9827e4d),
	.w8(32'h3bf2adab),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd4d2ee),
	.w1(32'h3b90d346),
	.w2(32'hba638f5a),
	.w3(32'hb9fee488),
	.w4(32'hbae027af),
	.w5(32'h3bbd226c),
	.w6(32'hbb1f7e4e),
	.w7(32'h3acc131a),
	.w8(32'h39f1f280),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0012c6),
	.w1(32'h3b3a0cda),
	.w2(32'hbb8b822c),
	.w3(32'h3b87ccde),
	.w4(32'hbb91b683),
	.w5(32'h3c294b1e),
	.w6(32'h3b4ea82b),
	.w7(32'hb87ad259),
	.w8(32'h3d298459),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39bb57cf),
	.w1(32'hbc4424e9),
	.w2(32'hbc878177),
	.w3(32'h3c505b2d),
	.w4(32'hbbaa43ae),
	.w5(32'h3a2d559e),
	.w6(32'h3c964366),
	.w7(32'hbc0f4f12),
	.w8(32'hbb02677a),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc00b34c),
	.w1(32'h3b55d137),
	.w2(32'hbbe96ab7),
	.w3(32'hb8260afe),
	.w4(32'hb8b908b2),
	.w5(32'hbc5fbaa2),
	.w6(32'h3b5148f9),
	.w7(32'h3ba3c0f3),
	.w8(32'hba8c9636),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbade8360),
	.w1(32'hb9c0c150),
	.w2(32'hba29c159),
	.w3(32'h3b1ea3ca),
	.w4(32'h3b4c3976),
	.w5(32'h3c026740),
	.w6(32'h3bf19b3e),
	.w7(32'h3ade6108),
	.w8(32'h3ba976ff),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae220c7),
	.w1(32'h3a84988f),
	.w2(32'h3af1441a),
	.w3(32'h3c16e638),
	.w4(32'h3c48ddba),
	.w5(32'h3a8b222a),
	.w6(32'h3c029a34),
	.w7(32'h3bb42659),
	.w8(32'h3a02e9c5),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d3f1e2),
	.w1(32'hbb08f754),
	.w2(32'h3afce132),
	.w3(32'hbadc260f),
	.w4(32'hbab80d98),
	.w5(32'hba2f1338),
	.w6(32'hbb9dea3c),
	.w7(32'h3ab9ea5a),
	.w8(32'h3b15e98d),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c176e55),
	.w1(32'h3a13cc67),
	.w2(32'h3aa1df66),
	.w3(32'hbb101edb),
	.w4(32'h3b1cfda5),
	.w5(32'h3c0e55ae),
	.w6(32'hbb364d5f),
	.w7(32'h3af3f649),
	.w8(32'h3b8dd596),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabf7f02),
	.w1(32'hba8fef90),
	.w2(32'hbb2c7835),
	.w3(32'h3ba33c00),
	.w4(32'hb89c0f15),
	.w5(32'hbbcbadfa),
	.w6(32'h3b4ea4b9),
	.w7(32'h3af9c5b8),
	.w8(32'hbb24cf57),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcad233),
	.w1(32'h3b336908),
	.w2(32'hba1ad6eb),
	.w3(32'h3ab36d64),
	.w4(32'hbab9485e),
	.w5(32'h3b4ab9ff),
	.w6(32'hbb94c6c7),
	.w7(32'hbb535aab),
	.w8(32'hbabd2661),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7a2332),
	.w1(32'hbb466cfd),
	.w2(32'hbc7d9c84),
	.w3(32'hbb8119cc),
	.w4(32'hbbc81d7c),
	.w5(32'hbc47805a),
	.w6(32'hbbe2c95f),
	.w7(32'hbb8993ad),
	.w8(32'hbbd24311),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2fcada),
	.w1(32'hbb7e1d8d),
	.w2(32'hbba9793f),
	.w3(32'hbc28350f),
	.w4(32'hbbc7d849),
	.w5(32'h3a8fcda2),
	.w6(32'hbbc92dd6),
	.w7(32'hbb2cd838),
	.w8(32'hbb12ffa8),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9b2e94),
	.w1(32'hbc5bf9c9),
	.w2(32'hbc0f533a),
	.w3(32'hbb71a0e5),
	.w4(32'hbb5fa368),
	.w5(32'hba071db1),
	.w6(32'hbb872397),
	.w7(32'hbb9571ab),
	.w8(32'h3aeeb2f1),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b50fbb1),
	.w1(32'hbb93b77f),
	.w2(32'hbc37a1a6),
	.w3(32'h3b41c3b9),
	.w4(32'h397baf59),
	.w5(32'hbc638a42),
	.w6(32'hbb37e3ba),
	.w7(32'hbbb981fb),
	.w8(32'hbc1e429c),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e866a3),
	.w1(32'h3b8dfb41),
	.w2(32'h3b85cb39),
	.w3(32'hbbe1d974),
	.w4(32'h3bd0259d),
	.w5(32'h3a09a9c9),
	.w6(32'hbae47499),
	.w7(32'h3bc5b56e),
	.w8(32'h3904a379),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be12f8e),
	.w1(32'h3bb05ddb),
	.w2(32'h39c7caa0),
	.w3(32'h3a2f605b),
	.w4(32'h3bd09592),
	.w5(32'hbae8d1fe),
	.w6(32'hba228d31),
	.w7(32'h3c420b85),
	.w8(32'h3b7f909c),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b517072),
	.w1(32'hbba97935),
	.w2(32'h3adf0b1b),
	.w3(32'hbbbe7cc6),
	.w4(32'hbb0aefba),
	.w5(32'hbbf24e81),
	.w6(32'hbbdf353e),
	.w7(32'h399c8c69),
	.w8(32'hbc1c0896),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd2e6b9),
	.w1(32'h3b0805b7),
	.w2(32'hbbed8899),
	.w3(32'h3b84101f),
	.w4(32'hbb98db43),
	.w5(32'hbb786300),
	.w6(32'hba86baed),
	.w7(32'hba5736e2),
	.w8(32'hbb37022e),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb78e660c),
	.w1(32'h3b828f64),
	.w2(32'h3c3abd26),
	.w3(32'hbb7899ee),
	.w4(32'h3c390e32),
	.w5(32'h3bbf15b7),
	.w6(32'hb9d74013),
	.w7(32'h3c460a49),
	.w8(32'h3b26c7c1),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab44486),
	.w1(32'hbb511784),
	.w2(32'hbb7566c1),
	.w3(32'hbb013adb),
	.w4(32'hbb3456ff),
	.w5(32'h3b01b99b),
	.w6(32'hbb604b81),
	.w7(32'h38771f09),
	.w8(32'h3a9b9a7d),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1fc2b7),
	.w1(32'hbb2030e0),
	.w2(32'h3aa870fc),
	.w3(32'hbaa73b96),
	.w4(32'h3aacbe4f),
	.w5(32'hbc17adff),
	.w6(32'hba089eb1),
	.w7(32'hba743d4f),
	.w8(32'hbc531a58),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc01ff60),
	.w1(32'h3b30c4a7),
	.w2(32'hbb566d30),
	.w3(32'hbc0af4c5),
	.w4(32'hbb33561d),
	.w5(32'hbc788078),
	.w6(32'hbb4bf2d7),
	.w7(32'h38d49108),
	.w8(32'hbc70e971),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0f8286),
	.w1(32'h3bed8a8d),
	.w2(32'h3b9a6d4b),
	.w3(32'hbb3fb4a2),
	.w4(32'hbab853a8),
	.w5(32'h3a537956),
	.w6(32'h3ba90aab),
	.w7(32'h3b3eb439),
	.w8(32'h39ad6870),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7ae8fb),
	.w1(32'hbc1c9446),
	.w2(32'hba6df540),
	.w3(32'hbb23382c),
	.w4(32'h3bcf23a0),
	.w5(32'hbbd36186),
	.w6(32'hbc1df607),
	.w7(32'h39679115),
	.w8(32'hbc458081),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399a4bb2),
	.w1(32'hbb2ca052),
	.w2(32'hbbce1cdc),
	.w3(32'hbba5e5ce),
	.w4(32'hbadb3824),
	.w5(32'h3b926c29),
	.w6(32'hbb7ae21a),
	.w7(32'h39b2c486),
	.w8(32'h3b5363ef),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9e2f453),
	.w1(32'hbb454593),
	.w2(32'hbbf56bbe),
	.w3(32'hbba44204),
	.w4(32'hbb8c35da),
	.w5(32'hba6059ef),
	.w6(32'hbbc41ac9),
	.w7(32'hbb2fcd99),
	.w8(32'h3ac32f8f),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb993f5e),
	.w1(32'hbbc6e821),
	.w2(32'hbbdba115),
	.w3(32'hba0bec10),
	.w4(32'hba3f32d3),
	.w5(32'h3bce26bb),
	.w6(32'hbb8aff54),
	.w7(32'hbbe903b2),
	.w8(32'h3bb243cb),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b307897),
	.w1(32'h3b4d1c2f),
	.w2(32'hbadffe4c),
	.w3(32'h3a465620),
	.w4(32'hb8c6f0ee),
	.w5(32'hbbe0f628),
	.w6(32'h3b10ba53),
	.w7(32'h3ae70b77),
	.w8(32'h3a23f655),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h384ebe61),
	.w1(32'hbb9118ac),
	.w2(32'hbc294f7c),
	.w3(32'hbbaefeec),
	.w4(32'hbaa877a4),
	.w5(32'h3b9ac9dd),
	.w6(32'h3c176efb),
	.w7(32'h3c0a59a8),
	.w8(32'h3c5f63aa),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h379048a2),
	.w1(32'hbb3e698c),
	.w2(32'hbba56f6e),
	.w3(32'hbb3f1cc4),
	.w4(32'hbc6ade00),
	.w5(32'h3b2d890d),
	.w6(32'hba7ed09c),
	.w7(32'hbc007d7d),
	.w8(32'h3bc244a9),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd37066),
	.w1(32'h3a828a7c),
	.w2(32'h3ad86a89),
	.w3(32'h3b19ae58),
	.w4(32'h3bad0c45),
	.w5(32'hb91c8401),
	.w6(32'h3b6ab679),
	.w7(32'h3b87278c),
	.w8(32'hbb5bfac9),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba041cb),
	.w1(32'h3a6d66b8),
	.w2(32'hba4011ed),
	.w3(32'h3a353651),
	.w4(32'hbb3e986a),
	.w5(32'hbc600b24),
	.w6(32'hbad26534),
	.w7(32'hbb292419),
	.w8(32'hbcaf22d2),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc82bb09),
	.w1(32'h3c46d7de),
	.w2(32'h3b32a126),
	.w3(32'hbc5940ef),
	.w4(32'hbc266d66),
	.w5(32'hbc13cd26),
	.w6(32'hbbb74823),
	.w7(32'hbacc6172),
	.w8(32'hbc5b0b22),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe90056),
	.w1(32'h398ab404),
	.w2(32'h3c162ad2),
	.w3(32'hbc3e9716),
	.w4(32'hbb45a89f),
	.w5(32'hbae159e4),
	.w6(32'hbb12b0b7),
	.w7(32'h3be0cfb7),
	.w8(32'hbb8118e7),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0a6d9f),
	.w1(32'hbbba24fe),
	.w2(32'hbc0b8130),
	.w3(32'hbb7c988c),
	.w4(32'hbbc4cf66),
	.w5(32'h3bb58e2b),
	.w6(32'hbc345b23),
	.w7(32'hbbdacb16),
	.w8(32'hbacab325),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9acf560),
	.w1(32'hbb617ec4),
	.w2(32'hbb9844c0),
	.w3(32'h3b27ed9f),
	.w4(32'hbb94820d),
	.w5(32'hbb42e7bd),
	.w6(32'hbc113c63),
	.w7(32'hbb8af11c),
	.w8(32'h3b10e36d),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc037416),
	.w1(32'hbb923fe3),
	.w2(32'hbb381004),
	.w3(32'hbbc18c13),
	.w4(32'hbbb2de4f),
	.w5(32'hbc8750aa),
	.w6(32'hbb724075),
	.w7(32'hbb09cdf6),
	.w8(32'hbc78665b),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad0b1f0),
	.w1(32'h3a031459),
	.w2(32'h3ba70b8f),
	.w3(32'hbbda8da9),
	.w4(32'h3b877302),
	.w5(32'h3bc12eda),
	.w6(32'hbc3ddccd),
	.w7(32'h3bb1c34f),
	.w8(32'hba4bc3c2),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb925b6d),
	.w1(32'h3b02697f),
	.w2(32'hbb69c987),
	.w3(32'h3be39682),
	.w4(32'hbb1a9209),
	.w5(32'hbb1421dc),
	.w6(32'h39c448e9),
	.w7(32'h3bc7a040),
	.w8(32'hbb47e703),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac95b8c),
	.w1(32'hb9de48e4),
	.w2(32'h3aadfe6b),
	.w3(32'hba9ca533),
	.w4(32'h3a0865b7),
	.w5(32'hbbc1670a),
	.w6(32'h3b0946b3),
	.w7(32'h3a9dd9c4),
	.w8(32'hb9bd1b40),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bca093b),
	.w1(32'hbbbd6572),
	.w2(32'hbc1c93a9),
	.w3(32'hbc151ab8),
	.w4(32'hb9b1a639),
	.w5(32'hbb13d913),
	.w6(32'hbbdc0868),
	.w7(32'hbba17be2),
	.w8(32'hbb28e511),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb920502),
	.w1(32'hbbd90a61),
	.w2(32'h39d25c76),
	.w3(32'hbb84194d),
	.w4(32'h3b2244dc),
	.w5(32'hbbc20ad6),
	.w6(32'hbc1e6378),
	.w7(32'h3ad46090),
	.w8(32'hbb3b3a09),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd7ebc2),
	.w1(32'hbc4b4539),
	.w2(32'hbb1e524c),
	.w3(32'hbbed58cd),
	.w4(32'hbc18cc1f),
	.w5(32'hbc16134d),
	.w6(32'h3b5b79b0),
	.w7(32'hbbe9b3dc),
	.w8(32'hbc08942d),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbce6e5),
	.w1(32'hbbaef2be),
	.w2(32'hbafaa983),
	.w3(32'hbb9c3416),
	.w4(32'h3b16c87f),
	.w5(32'hbc823d6d),
	.w6(32'hbc386ee3),
	.w7(32'h3b9698f3),
	.w8(32'hbc05114a),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf90224),
	.w1(32'hbc1ae2c7),
	.w2(32'hbc9abd81),
	.w3(32'hbc33dc52),
	.w4(32'hbbc005ab),
	.w5(32'h3c35974a),
	.w6(32'hbc14b21b),
	.w7(32'hbc733648),
	.w8(32'h3ca72347),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c7f43a2),
	.w1(32'h3c4849d9),
	.w2(32'hbc1211cb),
	.w3(32'h3c98cd91),
	.w4(32'h3bbef09d),
	.w5(32'hbb3f30cd),
	.w6(32'h3ce22aad),
	.w7(32'hbab167e0),
	.w8(32'hbb3a19a7),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3bbfdc),
	.w1(32'h3b1dcf08),
	.w2(32'hbb95ca6f),
	.w3(32'hbb8554c8),
	.w4(32'hbb958ce2),
	.w5(32'hbb4993bd),
	.w6(32'h380d1b0f),
	.w7(32'h3ac5165c),
	.w8(32'hbb41788a),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac6ec9e),
	.w1(32'hbb3f3e9a),
	.w2(32'hbb2df47c),
	.w3(32'hbc14b0fd),
	.w4(32'h3bb64ea3),
	.w5(32'h3a7ce51d),
	.w6(32'hbb6cf4f3),
	.w7(32'hbb4a299d),
	.w8(32'h3abce99c),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b425107),
	.w1(32'hbb58a676),
	.w2(32'hbb5330c9),
	.w3(32'h3b396ad8),
	.w4(32'hbbd5b2d4),
	.w5(32'hbbe9122d),
	.w6(32'hba0565e6),
	.w7(32'hbbd1f579),
	.w8(32'h3b2ffa00),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae57436),
	.w1(32'h3c25489f),
	.w2(32'hbbd0ae56),
	.w3(32'h3c4d3f07),
	.w4(32'h3a120f53),
	.w5(32'h3ab585e8),
	.w6(32'h3cd382c1),
	.w7(32'h3b7dc381),
	.w8(32'h3b99064b),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3371e9),
	.w1(32'h3b8b2855),
	.w2(32'hbb3e721c),
	.w3(32'h3a044f9a),
	.w4(32'hbb1e7d96),
	.w5(32'hbb2e57dc),
	.w6(32'h3bb150f6),
	.w7(32'hbbf44ef5),
	.w8(32'hbbd0f306),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8a6a65),
	.w1(32'hbb8fc533),
	.w2(32'h3899ca25),
	.w3(32'hba70311b),
	.w4(32'h3a93c755),
	.w5(32'h3965f5e9),
	.w6(32'hbbf21d9d),
	.w7(32'hbb748764),
	.w8(32'h392faf12),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b209825),
	.w1(32'hbb442981),
	.w2(32'h3ba1c10b),
	.w3(32'hba5da215),
	.w4(32'h3bbc5200),
	.w5(32'h3aee171d),
	.w6(32'hbbd3060c),
	.w7(32'h39f8309a),
	.w8(32'h3adb7e54),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b10cb3d),
	.w1(32'h3a79f6e8),
	.w2(32'h3acc3bea),
	.w3(32'hba241796),
	.w4(32'hba8d9569),
	.w5(32'h3c12ee2b),
	.w6(32'hba398cfb),
	.w7(32'h3abf69e1),
	.w8(32'h38d0c804),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4a4449),
	.w1(32'hbc9edfe7),
	.w2(32'h3c2f56b4),
	.w3(32'hbcb02ec3),
	.w4(32'h3a8313bd),
	.w5(32'hbbeb5996),
	.w6(32'hbc50848c),
	.w7(32'hbb67604e),
	.w8(32'hbb8df44a),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb777c09),
	.w1(32'hbb9010f8),
	.w2(32'h397ec1ee),
	.w3(32'hb9c88d3d),
	.w4(32'hb99791cd),
	.w5(32'h3b94ce54),
	.w6(32'hbb0778d6),
	.w7(32'hbb2b6981),
	.w8(32'h3c710ad6),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c2f637d),
	.w1(32'h3bbf6aab),
	.w2(32'h3b934a25),
	.w3(32'h3b9b4620),
	.w4(32'h3c9ad33f),
	.w5(32'hbc1b9a24),
	.w6(32'h3c38c292),
	.w7(32'h3d14323f),
	.w8(32'hbbdee29c),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6624e5),
	.w1(32'h39490c78),
	.w2(32'h3b801ab6),
	.w3(32'hbaedaa10),
	.w4(32'h3c0340e2),
	.w5(32'h3be43585),
	.w6(32'hbc20babd),
	.w7(32'h3ac20147),
	.w8(32'h3b88eac5),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3c9d3e),
	.w1(32'hbc5408cd),
	.w2(32'hba70cb30),
	.w3(32'hbc21b27d),
	.w4(32'hbbc86c9a),
	.w5(32'hba5f5714),
	.w6(32'hbc101b6f),
	.w7(32'hbc0653e6),
	.w8(32'hba930211),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb29a8d8),
	.w1(32'hbaa5ca31),
	.w2(32'h3ad12a05),
	.w3(32'hbb1668b9),
	.w4(32'h3aa14bc5),
	.w5(32'h380e94b3),
	.w6(32'hbb874125),
	.w7(32'hba0c16bd),
	.w8(32'hbaa1c501),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a683a6e),
	.w1(32'hbc3f10c6),
	.w2(32'hbb55a19f),
	.w3(32'hbbfea654),
	.w4(32'hbc1ff0f2),
	.w5(32'hbb6f1dae),
	.w6(32'hba6b4a6f),
	.w7(32'hbc011d55),
	.w8(32'h3a456393),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba30f2c),
	.w1(32'hbbbed10c),
	.w2(32'hba7517e3),
	.w3(32'h3b4c5b23),
	.w4(32'h3b9a5f45),
	.w5(32'hba9c8ecc),
	.w6(32'h3ae28f64),
	.w7(32'h39aa1b6b),
	.w8(32'h3a92551c),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb428425),
	.w1(32'h3abb5005),
	.w2(32'hbc0a2679),
	.w3(32'h3be7de87),
	.w4(32'hbb943500),
	.w5(32'h3c6e1f87),
	.w6(32'h3c1c8972),
	.w7(32'hbb779fd0),
	.w8(32'h3c3fd7ec),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ce34ad6),
	.w1(32'hbbdb2fb5),
	.w2(32'h3c8357ab),
	.w3(32'hbc4551ab),
	.w4(32'h39fd67f5),
	.w5(32'hbb0dddae),
	.w6(32'hbbd3e5c8),
	.w7(32'hbc1fd1f8),
	.w8(32'h3b719859),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b91bc53),
	.w1(32'h3c344927),
	.w2(32'h3af434a9),
	.w3(32'hba1a1be6),
	.w4(32'h3b2fbf64),
	.w5(32'h3b77f876),
	.w6(32'h3c8fce72),
	.w7(32'h3a9d248e),
	.w8(32'hbae3c5b3),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba13e182),
	.w1(32'hbc019ee4),
	.w2(32'hbbfb50d4),
	.w3(32'hbba6c894),
	.w4(32'hbbb8a82a),
	.w5(32'h3a6dd8ff),
	.w6(32'hbbb8aaa9),
	.w7(32'hba29f0db),
	.w8(32'h3b476378),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af123b5),
	.w1(32'h3b5944e7),
	.w2(32'hbb9d3750),
	.w3(32'hbb6933f5),
	.w4(32'hbb477ed2),
	.w5(32'h3b0e9a13),
	.w6(32'hbb935b6b),
	.w7(32'hbb2d5896),
	.w8(32'h3b1ca1c1),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8b65fa),
	.w1(32'hbaa738f1),
	.w2(32'hbb69a1ae),
	.w3(32'h3a9e71ab),
	.w4(32'hb97c42cd),
	.w5(32'h3c40ef68),
	.w6(32'h3ac5a191),
	.w7(32'h3b78dd7c),
	.w8(32'h3bf23aca),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be7aa57),
	.w1(32'hbc2c6b53),
	.w2(32'h3ba28080),
	.w3(32'hbc526a0c),
	.w4(32'h3c50b0fe),
	.w5(32'hbb46cd3c),
	.w6(32'hbc7cf60d),
	.w7(32'hbb194372),
	.w8(32'hbb21de3f),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd6fcc1),
	.w1(32'hba075d09),
	.w2(32'h383500e6),
	.w3(32'hba88667c),
	.w4(32'hb9b19a3f),
	.w5(32'h3b91f469),
	.w6(32'hbb5a931e),
	.w7(32'hbb86bf0d),
	.w8(32'h3be7e72d),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba522b2b),
	.w1(32'h3b265ac6),
	.w2(32'h3c33e8a6),
	.w3(32'hbbb43f15),
	.w4(32'h3c0b48d3),
	.w5(32'hba4963c5),
	.w6(32'hbbd9bd24),
	.w7(32'h3bf8cf7b),
	.w8(32'hb9c80418),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule