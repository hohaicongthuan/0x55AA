module layer_10_featuremap_327(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39d3e6c3),
	.w1(32'hb998fbbb),
	.w2(32'h3a975538),
	.w3(32'h3a8ae315),
	.w4(32'h3ad32ede),
	.w5(32'h39096119),
	.w6(32'h39f2f7cb),
	.w7(32'h3a969a8d),
	.w8(32'h39bdef71),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb984ed27),
	.w1(32'hb94ec784),
	.w2(32'h3a171ea0),
	.w3(32'hb91f676c),
	.w4(32'h3a452294),
	.w5(32'h3a0dfbf4),
	.w6(32'h37cfdf0c),
	.w7(32'h397d2c67),
	.w8(32'hb9ad4076),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba84fcb3),
	.w1(32'h391bc0fd),
	.w2(32'h394120e8),
	.w3(32'hb9b03ad2),
	.w4(32'h384a2e14),
	.w5(32'h399aec36),
	.w6(32'hb9af2275),
	.w7(32'hb796315f),
	.w8(32'h39f3f738),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2d55fc),
	.w1(32'h3a593314),
	.w2(32'h3aa843fc),
	.w3(32'h38e958c3),
	.w4(32'h3a3b16c8),
	.w5(32'hba5ec5fd),
	.w6(32'h38b8bd49),
	.w7(32'h3a7e5116),
	.w8(32'hbabb2149),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ed2c8f),
	.w1(32'hba90e261),
	.w2(32'hba8e0074),
	.w3(32'hbab88373),
	.w4(32'hba320ea6),
	.w5(32'h39a9a446),
	.w6(32'hbb29a629),
	.w7(32'hbae15798),
	.w8(32'h38acbbac),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b10294),
	.w1(32'hb98a4a48),
	.w2(32'h39fa0691),
	.w3(32'hb8dfdfdb),
	.w4(32'h3a57ba92),
	.w5(32'h39916b65),
	.w6(32'hba091023),
	.w7(32'h39b75900),
	.w8(32'h39a20778),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aae0543),
	.w1(32'hb9497165),
	.w2(32'hba9bff60),
	.w3(32'h385a923a),
	.w4(32'hb98371ee),
	.w5(32'hba384d18),
	.w6(32'h3a103c37),
	.w7(32'hba0a9a15),
	.w8(32'hba8213bf),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98ab00a),
	.w1(32'hbabcba75),
	.w2(32'h3998f2c9),
	.w3(32'hbad76d14),
	.w4(32'hb9c11996),
	.w5(32'h3a5c63d2),
	.w6(32'hbaf75861),
	.w7(32'hb9442e0c),
	.w8(32'h388358e8),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6a9df0),
	.w1(32'h3a18cc54),
	.w2(32'h3a82dceb),
	.w3(32'h3a390081),
	.w4(32'h3ad40e66),
	.w5(32'h3a140c27),
	.w6(32'h3a1be624),
	.w7(32'h3a822fbe),
	.w8(32'h39995695),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a078de6),
	.w1(32'h39a074b2),
	.w2(32'h39c5aa81),
	.w3(32'h384ef7d4),
	.w4(32'h3a992096),
	.w5(32'h391918c7),
	.w6(32'hba3caad4),
	.w7(32'hb750364a),
	.w8(32'hba462508),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f09a3e),
	.w1(32'h386fad66),
	.w2(32'h3a749a6a),
	.w3(32'h38878e30),
	.w4(32'h3a5000e7),
	.w5(32'h391612ec),
	.w6(32'hb89d0f90),
	.w7(32'h3a3a2886),
	.w8(32'h39e56b87),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a93f60d),
	.w1(32'h3aa90714),
	.w2(32'hba125eb9),
	.w3(32'h382baffc),
	.w4(32'hb9c1e9e9),
	.w5(32'hbb1ded6e),
	.w6(32'h39cef189),
	.w7(32'h38097a5e),
	.w8(32'hbafc4de7),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9cbf4b3),
	.w1(32'hba185144),
	.w2(32'hbacedfa2),
	.w3(32'hb97c5d22),
	.w4(32'hba66d950),
	.w5(32'hba075b60),
	.w6(32'hba0772e9),
	.w7(32'hbac39b71),
	.w8(32'hbab237be),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8f9485c),
	.w1(32'hba74160e),
	.w2(32'hb78c7311),
	.w3(32'hb9ff2f46),
	.w4(32'hb928df8a),
	.w5(32'hba0c9777),
	.w6(32'hb98bd6d2),
	.w7(32'hb9c4209e),
	.w8(32'hb9c71fe5),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f88552),
	.w1(32'h3916f8e8),
	.w2(32'h388685c4),
	.w3(32'hba0fc66d),
	.w4(32'h3a8904fc),
	.w5(32'h384a505a),
	.w6(32'hba2cc897),
	.w7(32'h3976de23),
	.w8(32'hb9b516fb),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9dd6a0f),
	.w1(32'hba4f8ead),
	.w2(32'hba69f27e),
	.w3(32'hb9bd349c),
	.w4(32'h39fd0084),
	.w5(32'h3a98128b),
	.w6(32'hba3d19ce),
	.w7(32'hb9e6d2a1),
	.w8(32'hba3182f3),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3886b989),
	.w1(32'hb9fb9f78),
	.w2(32'h394eeaf7),
	.w3(32'h3a527c8b),
	.w4(32'h3a61215d),
	.w5(32'hb981ed83),
	.w6(32'h370c814e),
	.w7(32'h39a6be60),
	.w8(32'hba2aa155),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a79450),
	.w1(32'hbac34356),
	.w2(32'hbafc1fcf),
	.w3(32'h36d5ba6b),
	.w4(32'hba6c432e),
	.w5(32'hbabc92d6),
	.w6(32'hbaa760da),
	.w7(32'hba9caebd),
	.w8(32'hbb05ee86),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39991d39),
	.w1(32'hbabc9f9e),
	.w2(32'hbae4f3bd),
	.w3(32'hb91fd4ca),
	.w4(32'hba96b292),
	.w5(32'hbaa23d42),
	.w6(32'hbaa78a11),
	.w7(32'hbaafb19e),
	.w8(32'hbaa6262e),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98b1620),
	.w1(32'hb7ac4066),
	.w2(32'hba1c65d1),
	.w3(32'hb9faa433),
	.w4(32'hb906e657),
	.w5(32'h39575b53),
	.w6(32'hb9601378),
	.w7(32'hba068443),
	.w8(32'h39832935),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a382d2d),
	.w1(32'h39b4f2a4),
	.w2(32'hb9450793),
	.w3(32'hb972904e),
	.w4(32'h390a9526),
	.w5(32'h3aa9f75e),
	.w6(32'h3a04fe6d),
	.w7(32'h394a9028),
	.w8(32'h3ab90acf),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab3d5de),
	.w1(32'h3ae01fba),
	.w2(32'h3aa9a1b0),
	.w3(32'h3a82c281),
	.w4(32'h3aa788ba),
	.w5(32'hb89a9bec),
	.w6(32'h3a29b0a6),
	.w7(32'h3a8fef19),
	.w8(32'hb98c78da),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb285442),
	.w1(32'hba879a55),
	.w2(32'hbb091aaf),
	.w3(32'hbae5e6e0),
	.w4(32'hba939bc3),
	.w5(32'hbac9b8e6),
	.w6(32'hbb175030),
	.w7(32'hbabc177f),
	.w8(32'hbb1e2893),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba23f497),
	.w1(32'hba11e796),
	.w2(32'hb967aed9),
	.w3(32'hbab75cb7),
	.w4(32'h38864982),
	.w5(32'h3a73885c),
	.w6(32'hbabcea71),
	.w7(32'hb9f91184),
	.w8(32'hba77a3bb),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb08142a),
	.w1(32'h3a2716a8),
	.w2(32'h39e6b1ae),
	.w3(32'hba7a5a19),
	.w4(32'h39f3f140),
	.w5(32'h3a8bebf1),
	.w6(32'hbb24aacd),
	.w7(32'h3972d3bc),
	.w8(32'hba68f823),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c14101),
	.w1(32'h3a3913b6),
	.w2(32'h3992e896),
	.w3(32'h3a54ea42),
	.w4(32'h3a41602d),
	.w5(32'hba1f4427),
	.w6(32'h3a69fb7e),
	.w7(32'h39b835f1),
	.w8(32'hba672700),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba93c338),
	.w1(32'hba87991e),
	.w2(32'hbacd52a5),
	.w3(32'hba5739ed),
	.w4(32'hbaa6cf0d),
	.w5(32'h3aae3ce0),
	.w6(32'hba2c0003),
	.w7(32'hbaaf8024),
	.w8(32'h3a7845c6),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b29f5cc),
	.w1(32'h38d4f236),
	.w2(32'h39b3a5b9),
	.w3(32'h3aafe9f8),
	.w4(32'h3ae4829a),
	.w5(32'hba1e0b9b),
	.w6(32'h3a454658),
	.w7(32'h3a5b8c41),
	.w8(32'hbad00089),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba94a660),
	.w1(32'hba5b2393),
	.w2(32'hb9b18932),
	.w3(32'hba52866b),
	.w4(32'hb9683391),
	.w5(32'hb7bd931b),
	.w6(32'hba8a2dd2),
	.w7(32'hba187aa3),
	.w8(32'hb9debaaf),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8e9a5e),
	.w1(32'h3989ff4a),
	.w2(32'h3a6fca93),
	.w3(32'h39cd1a33),
	.w4(32'h3a829034),
	.w5(32'hb8e3314b),
	.w6(32'h398816fc),
	.w7(32'h3a028678),
	.w8(32'hba74b407),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b4f0ce),
	.w1(32'hb9d54847),
	.w2(32'hba412a70),
	.w3(32'hbac53222),
	.w4(32'hb9b7e0d8),
	.w5(32'h394f7a69),
	.w6(32'hba57d997),
	.w7(32'h3940038a),
	.w8(32'h39fb065c),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8c2cf98),
	.w1(32'hb9edd886),
	.w2(32'hb8a6931e),
	.w3(32'h39c729c7),
	.w4(32'h38f0d532),
	.w5(32'h3978e1f9),
	.w6(32'h394405a1),
	.w7(32'h39e56a72),
	.w8(32'h3989e02b),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a76d0c3),
	.w1(32'h393c9111),
	.w2(32'h38b2c66d),
	.w3(32'h3a363588),
	.w4(32'h3a54a338),
	.w5(32'hb9ab7be1),
	.w6(32'h39ff6e23),
	.w7(32'h3a08b72f),
	.w8(32'hba768cc2),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9c37af),
	.w1(32'hb9f0e044),
	.w2(32'h38f69d40),
	.w3(32'hba6930b1),
	.w4(32'h39bd93a1),
	.w5(32'hb8ef2c0f),
	.w6(32'hba99732a),
	.w7(32'hb87b13b1),
	.w8(32'hb94d1446),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39b2b641),
	.w1(32'hb8d8f256),
	.w2(32'h388a47bb),
	.w3(32'h39314b61),
	.w4(32'h3934447b),
	.w5(32'h3a364de6),
	.w6(32'h389aef54),
	.w7(32'hb889ece6),
	.w8(32'hba52f816),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3906ef07),
	.w1(32'hb7e3f027),
	.w2(32'h392129e4),
	.w3(32'hb791a944),
	.w4(32'hb7e6663b),
	.w5(32'hb9297ae5),
	.w6(32'hba320528),
	.w7(32'hb8c96bd9),
	.w8(32'hb8f1472b),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac87f7e),
	.w1(32'h3aba6432),
	.w2(32'hbb1e27e9),
	.w3(32'hb9e9cb68),
	.w4(32'h3b01b264),
	.w5(32'hb9be50d0),
	.w6(32'hba8d2d15),
	.w7(32'h3a61b901),
	.w8(32'hba5c6efb),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadf492a),
	.w1(32'h3a786261),
	.w2(32'hb8ac5c79),
	.w3(32'hb7583406),
	.w4(32'h3b2159cf),
	.w5(32'h3a9a7833),
	.w6(32'hbade9ec3),
	.w7(32'h3a36e29a),
	.w8(32'hba1c19af),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9a9122),
	.w1(32'h3894271a),
	.w2(32'h37f8f935),
	.w3(32'hba44fe31),
	.w4(32'h3992586b),
	.w5(32'h399d2959),
	.w6(32'hbaacef50),
	.w7(32'hb98f685e),
	.w8(32'hba42c501),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39355125),
	.w1(32'h39e3ff8b),
	.w2(32'h3a6cb05a),
	.w3(32'h3a5a9467),
	.w4(32'h3ae86b83),
	.w5(32'h390c6012),
	.w6(32'hb99e1ad5),
	.w7(32'h3a874516),
	.w8(32'hb9d3cfc0),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9d9b38e),
	.w1(32'hba0aa6df),
	.w2(32'h3957e6ab),
	.w3(32'hb99354c8),
	.w4(32'hb9323f5b),
	.w5(32'h3a65b966),
	.w6(32'h3950adf5),
	.w7(32'hb9974cc6),
	.w8(32'h39a300f1),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a128a69),
	.w1(32'h3a5a04dd),
	.w2(32'h3a4e8d41),
	.w3(32'h3a686c40),
	.w4(32'h3a36761b),
	.w5(32'h39be759e),
	.w6(32'h3a757c4a),
	.w7(32'h39ba5b58),
	.w8(32'hba0efcc1),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0406bd),
	.w1(32'hba4233cc),
	.w2(32'hb950281c),
	.w3(32'hb88906be),
	.w4(32'h3a07c07b),
	.w5(32'hba99a625),
	.w6(32'hba866a54),
	.w7(32'hb91f5066),
	.w8(32'hbaf76f61),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac5d6c0),
	.w1(32'hbb392efe),
	.w2(32'hbb0ca0fd),
	.w3(32'hbac0adef),
	.w4(32'hbac2dc9e),
	.w5(32'hba3b40e0),
	.w6(32'hbb2a542b),
	.w7(32'hbb2e1783),
	.w8(32'hbaea83f5),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab25fc2),
	.w1(32'hba071a5b),
	.w2(32'hb9eb50ae),
	.w3(32'hba800212),
	.w4(32'h399e042c),
	.w5(32'hba182a4b),
	.w6(32'hbb090416),
	.w7(32'hba4d0a20),
	.w8(32'hbb01367a),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf8e3e5),
	.w1(32'h3853603f),
	.w2(32'hb9593e64),
	.w3(32'hbaba690d),
	.w4(32'h3944c95c),
	.w5(32'hba219f01),
	.w6(32'hbb25a3ca),
	.w7(32'hba5a8d52),
	.w8(32'hbb0b5f11),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba86f685),
	.w1(32'hb950f463),
	.w2(32'hba1ffed9),
	.w3(32'hbab7d920),
	.w4(32'hb938ee11),
	.w5(32'h3b1a4925),
	.w6(32'hbb0dfd1f),
	.w7(32'hba86060b),
	.w8(32'h3aba873c),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b668c10),
	.w1(32'h3ad5990f),
	.w2(32'h386e5bcd),
	.w3(32'h3b2492e0),
	.w4(32'h3a9ca550),
	.w5(32'hbb2c011f),
	.w6(32'h3a9e33b3),
	.w7(32'h39831bd5),
	.w8(32'hbb55d4b4),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba678575),
	.w1(32'hba100c52),
	.w2(32'hb98824c8),
	.w3(32'hba171e17),
	.w4(32'h37424a70),
	.w5(32'h3ae0e3d0),
	.w6(32'hba0b2622),
	.w7(32'hb9c75d69),
	.w8(32'h3af34446),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aece5ff),
	.w1(32'h3aea2930),
	.w2(32'h3ad3b0ad),
	.w3(32'h3aaae3ef),
	.w4(32'h3ac2f0e1),
	.w5(32'hba1697c4),
	.w6(32'h3aa49bbc),
	.w7(32'h3a8b0351),
	.w8(32'hb9a2acee),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a22d306),
	.w1(32'hba5ade22),
	.w2(32'hba6dc9c4),
	.w3(32'hba602a4b),
	.w4(32'hb99ae45b),
	.w5(32'h393d1adf),
	.w6(32'hbac71ad6),
	.w7(32'hba8d0c25),
	.w8(32'h3a398fed),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa2d8fe),
	.w1(32'hba7fdf43),
	.w2(32'hb940e7cf),
	.w3(32'hba48d3a7),
	.w4(32'hb9d45f64),
	.w5(32'hb85a9b5e),
	.w6(32'hbaa1f17f),
	.w7(32'hb764246d),
	.w8(32'hba6ff301),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb99877d3),
	.w1(32'hba323d64),
	.w2(32'hb806cb8b),
	.w3(32'hba149d25),
	.w4(32'hba51591e),
	.w5(32'h39bfc2c0),
	.w6(32'hba5bb909),
	.w7(32'hba544c33),
	.w8(32'h3a345ebd),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa12daf),
	.w1(32'hba00cf10),
	.w2(32'hbaeea43e),
	.w3(32'h387e9a06),
	.w4(32'hb928a454),
	.w5(32'hbaec72b3),
	.w6(32'h385e63e4),
	.w7(32'hbaea6e97),
	.w8(32'hbabda5b0),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7d67975),
	.w1(32'hba0911bb),
	.w2(32'hba80be14),
	.w3(32'hb993be9c),
	.w4(32'h39746ecf),
	.w5(32'hba19158b),
	.w6(32'hb9decff7),
	.w7(32'hb9dbe94b),
	.w8(32'hba2da561),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb90293dd),
	.w1(32'hba30000d),
	.w2(32'h38a8a36f),
	.w3(32'h38b1d41c),
	.w4(32'h39e5a599),
	.w5(32'h38f622f2),
	.w6(32'hb9b83917),
	.w7(32'hb8c23524),
	.w8(32'h387892fa),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h399262d3),
	.w1(32'h392551aa),
	.w2(32'h39765ad8),
	.w3(32'h3947e3cc),
	.w4(32'h3995a5f1),
	.w5(32'hba721ebe),
	.w6(32'h39ce2609),
	.w7(32'h38a0655e),
	.w8(32'hba5730fb),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4cf7ae),
	.w1(32'hba70653a),
	.w2(32'hba316598),
	.w3(32'hbabd53cd),
	.w4(32'hb9ecf019),
	.w5(32'h3af11aed),
	.w6(32'hbab608fa),
	.w7(32'hba8b3749),
	.w8(32'h3af1a2f6),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aff5e0f),
	.w1(32'h3af8a89e),
	.w2(32'h3ae0e873),
	.w3(32'h3acec018),
	.w4(32'h3aef18fa),
	.w5(32'h3a0d3e5e),
	.w6(32'h3ad8359e),
	.w7(32'h3aacb993),
	.w8(32'hba2caae6),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a51b736),
	.w1(32'h3a3e64ee),
	.w2(32'h3a61d640),
	.w3(32'h39c3ad2f),
	.w4(32'h3975fdaf),
	.w5(32'hb95aa34d),
	.w6(32'hbade0cb8),
	.w7(32'hba2dd258),
	.w8(32'h38cefac5),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3948ab19),
	.w1(32'h383b92d2),
	.w2(32'hb9f3d19b),
	.w3(32'hb95c20c2),
	.w4(32'h38787fd4),
	.w5(32'h3988a8fa),
	.w6(32'hba07f27f),
	.w7(32'hb9e1a7f1),
	.w8(32'hb90325e1),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394405bb),
	.w1(32'hb8bbc449),
	.w2(32'hb924a631),
	.w3(32'h3a1bb8d0),
	.w4(32'h392e372a),
	.w5(32'hba999ad1),
	.w6(32'h39c12b9b),
	.w7(32'h39b846a8),
	.w8(32'hbaab73ed),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9f63172),
	.w1(32'hba2ae8da),
	.w2(32'hba056063),
	.w3(32'hba77de51),
	.w4(32'hb9c62d27),
	.w5(32'hb9dfe357),
	.w6(32'hba9e566a),
	.w7(32'hb9bd4b1e),
	.w8(32'hba3d38f8),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba106b05),
	.w1(32'hba5b6454),
	.w2(32'hb970c6bc),
	.w3(32'hba28f905),
	.w4(32'hb95dd1ff),
	.w5(32'hb8dbbc8a),
	.w6(32'hb989626d),
	.w7(32'hba58481f),
	.w8(32'h39db4000),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0f0356),
	.w1(32'hb9c04829),
	.w2(32'hba7e46f8),
	.w3(32'hb9563d11),
	.w4(32'h394a9767),
	.w5(32'hb9b0a3b7),
	.w6(32'hb9fbe2d8),
	.w7(32'hba4aec15),
	.w8(32'hb9d621d4),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7b0fe3e),
	.w1(32'hb9fa272d),
	.w2(32'hb9b3408b),
	.w3(32'hb984b7d1),
	.w4(32'h39d135e0),
	.w5(32'h3a1434aa),
	.w6(32'hbaa7a651),
	.w7(32'hb8823e58),
	.w8(32'h3a13cfec),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a90b57f),
	.w1(32'hb98b8c5e),
	.w2(32'h39463ac5),
	.w3(32'h3a60d03e),
	.w4(32'h3a07972c),
	.w5(32'hbb06cd2e),
	.w6(32'h3947da59),
	.w7(32'h39cb8bb7),
	.w8(32'hbb4f4ed8),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf8c463),
	.w1(32'hba38dc62),
	.w2(32'hba49b8b6),
	.w3(32'hbac176ce),
	.w4(32'hba5097af),
	.w5(32'h3846b5ee),
	.w6(32'hbad581f0),
	.w7(32'hbae1a246),
	.w8(32'hbaa3d82a),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9afa6fd),
	.w1(32'hba24af72),
	.w2(32'hba9cbdb8),
	.w3(32'hba2976f0),
	.w4(32'hb9cc86dc),
	.w5(32'hba54b076),
	.w6(32'hba530f73),
	.w7(32'hbaa0677e),
	.w8(32'hbb39e1e8),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2726d5),
	.w1(32'hba5a5961),
	.w2(32'hba0b1746),
	.w3(32'hbabef2aa),
	.w4(32'h3ac8394b),
	.w5(32'h39a784f8),
	.w6(32'hbb8776e3),
	.w7(32'hba94f30c),
	.w8(32'hbad0a527),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c29bdc),
	.w1(32'hba9e7bdf),
	.w2(32'hba3ed63e),
	.w3(32'hb9d703e9),
	.w4(32'hba3d456a),
	.w5(32'h3a438f6b),
	.w6(32'hbab52feb),
	.w7(32'hba559a7e),
	.w8(32'h360120fb),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3988e722),
	.w1(32'h387f7f2e),
	.w2(32'hb97ebc44),
	.w3(32'h38335977),
	.w4(32'hba6079ba),
	.w5(32'h3a929127),
	.w6(32'h371868bb),
	.w7(32'h38e7c62b),
	.w8(32'h393c7845),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1b8e97),
	.w1(32'h3a9ad5eb),
	.w2(32'h3a33d7bc),
	.w3(32'h3a969d13),
	.w4(32'h3a5d3305),
	.w5(32'hb99080f4),
	.w6(32'h3a6b1986),
	.w7(32'h3a8088fa),
	.w8(32'hb9cbef14),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a9a38a),
	.w1(32'hba0dc2cb),
	.w2(32'hba9675b6),
	.w3(32'h380807f8),
	.w4(32'hba3f2d16),
	.w5(32'h398cb9e9),
	.w6(32'hb921aadc),
	.w7(32'hba84073d),
	.w8(32'h39816acd),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h374e879f),
	.w1(32'hb9d26674),
	.w2(32'h3a7a9376),
	.w3(32'h38a5a59d),
	.w4(32'h3a8267c1),
	.w5(32'hba692a57),
	.w6(32'h38015502),
	.w7(32'h3a4bce01),
	.w8(32'hbab8d5f9),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9abe29c),
	.w1(32'hba622a04),
	.w2(32'hbadae649),
	.w3(32'hba094533),
	.w4(32'hba400df0),
	.w5(32'hba8e0101),
	.w6(32'hbaa0cf39),
	.w7(32'hbae586b0),
	.w8(32'hba88f053),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38b2ec6d),
	.w1(32'hb9902142),
	.w2(32'hba78e76c),
	.w3(32'hba4f08c4),
	.w4(32'h39f0e58d),
	.w5(32'hbb038c05),
	.w6(32'hbadd57af),
	.w7(32'hba653246),
	.w8(32'hbad7ca81),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9d5211),
	.w1(32'hbaae6096),
	.w2(32'hb9a62dde),
	.w3(32'hba8760f5),
	.w4(32'h396a8514),
	.w5(32'hba8c5eed),
	.w6(32'hbb264997),
	.w7(32'hba0ad848),
	.w8(32'hbb0425d5),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabbe9a6),
	.w1(32'hbad31681),
	.w2(32'hbacfb4da),
	.w3(32'hbad45426),
	.w4(32'hbaaf32d3),
	.w5(32'hb824d25f),
	.w6(32'hbb1f1d30),
	.w7(32'hbab62de4),
	.w8(32'hba4d6f71),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7e2a18),
	.w1(32'hb7c20b2b),
	.w2(32'h39a5f9df),
	.w3(32'h37dbedd9),
	.w4(32'h3a7af645),
	.w5(32'hb7002c78),
	.w6(32'hb8d4c047),
	.w7(32'h39d80d4a),
	.w8(32'hb99f4b03),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba388b0a),
	.w1(32'h38c81ac1),
	.w2(32'hb9cac9e8),
	.w3(32'hba0a9927),
	.w4(32'hb8ebfee0),
	.w5(32'h3a18585e),
	.w6(32'h38c54767),
	.w7(32'hb6fbde69),
	.w8(32'hba21d451),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39c4e18d),
	.w1(32'hba159ae0),
	.w2(32'hba7c7ad1),
	.w3(32'h3a316028),
	.w4(32'h39888d16),
	.w5(32'hb88a9b6c),
	.w6(32'hba27d2a2),
	.w7(32'hba1b3c26),
	.w8(32'hb9cc9457),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39430b51),
	.w1(32'h39979867),
	.w2(32'h39edfd23),
	.w3(32'h3820c292),
	.w4(32'h37c0a614),
	.w5(32'hba2e55af),
	.w6(32'hb8d4707a),
	.w7(32'hb7630a9a),
	.w8(32'hba79f27f),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba879b48),
	.w1(32'h37c8f7ec),
	.w2(32'hb83ef718),
	.w3(32'hb9306685),
	.w4(32'hb950151c),
	.w5(32'h3912abfe),
	.w6(32'h3a6acb75),
	.w7(32'h39bdba40),
	.w8(32'hb9e01ec5),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2ea1f0),
	.w1(32'hb9b8ca54),
	.w2(32'h38825dba),
	.w3(32'hb873ddff),
	.w4(32'hb9c38c6f),
	.w5(32'hb9221d49),
	.w6(32'hb9f20405),
	.w7(32'hb96ebe65),
	.w8(32'hba80f7a2),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5d1d49),
	.w1(32'h39b09c5c),
	.w2(32'h39bd0ae9),
	.w3(32'h38a05af5),
	.w4(32'h39a6308b),
	.w5(32'h39907df0),
	.w6(32'hb9511c07),
	.w7(32'h399fa9d6),
	.w8(32'h39e8fd17),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba820ca2),
	.w1(32'h39e9ee32),
	.w2(32'hba060a3b),
	.w3(32'hbaa7cb1a),
	.w4(32'h3aa82a51),
	.w5(32'hb7ef89ba),
	.w6(32'hba51572b),
	.w7(32'hb9095f95),
	.w8(32'hba529cc5),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9baf267),
	.w1(32'hb95043c4),
	.w2(32'hb9229392),
	.w3(32'hb9c532fa),
	.w4(32'hb9824fb7),
	.w5(32'h39de408f),
	.w6(32'hba4c6c15),
	.w7(32'hb8b5ae71),
	.w8(32'h39c6b2eb),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3787e331),
	.w1(32'hb88d4f5b),
	.w2(32'hb6ee423d),
	.w3(32'hb8f5ead5),
	.w4(32'h3a669321),
	.w5(32'h391fd6c1),
	.w6(32'hba10d5a1),
	.w7(32'hb698302e),
	.w8(32'hba49adf9),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba5ab2ec),
	.w1(32'hb93461fb),
	.w2(32'h3a8e17b8),
	.w3(32'hb80370ef),
	.w4(32'h3a90868b),
	.w5(32'hbb0a34fa),
	.w6(32'h389d2ff6),
	.w7(32'h39b7ee02),
	.w8(32'hbadee10a),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7ae526),
	.w1(32'hba4ad08c),
	.w2(32'hb8e48a99),
	.w3(32'hba6262ea),
	.w4(32'h390c61f4),
	.w5(32'hbb0d9534),
	.w6(32'hba157abf),
	.w7(32'hb91c9460),
	.w8(32'hbb1e16ad),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad5dc4e),
	.w1(32'h3a6a6971),
	.w2(32'h3a2c89fa),
	.w3(32'h3a3c667e),
	.w4(32'h3ac57f5a),
	.w5(32'hbac92f5c),
	.w6(32'h3a0a1ea1),
	.w7(32'h3a8e4d51),
	.w8(32'hbb0e2d48),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb00382e),
	.w1(32'hbb1bebfc),
	.w2(32'hba9c68b7),
	.w3(32'hba52926b),
	.w4(32'hb8d0ba48),
	.w5(32'hba581ac1),
	.w6(32'hba792ea1),
	.w7(32'hba98037b),
	.w8(32'hba9ace17),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba418f91),
	.w1(32'hbaa63676),
	.w2(32'hb88eb1b3),
	.w3(32'hbaa32db9),
	.w4(32'h39c8b079),
	.w5(32'h39d97c0a),
	.w6(32'hbaf8ab3f),
	.w7(32'h382d5749),
	.w8(32'hba8b9c3c),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba739033),
	.w1(32'hb940a4a4),
	.w2(32'h38cda6e1),
	.w3(32'h39797816),
	.w4(32'h39fb3fdc),
	.w5(32'h398b1d99),
	.w6(32'h3663e94c),
	.w7(32'h397e7df6),
	.w8(32'hb95dff93),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9b6984),
	.w1(32'h38a7859e),
	.w2(32'hb9ebb65c),
	.w3(32'hba1d873a),
	.w4(32'h3a6fb3be),
	.w5(32'hba18e70e),
	.w6(32'hbac6a46a),
	.w7(32'hba03dc11),
	.w8(32'hbacc3988),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8a8e26),
	.w1(32'hba789240),
	.w2(32'hbad05d2c),
	.w3(32'hba867949),
	.w4(32'hbacad183),
	.w5(32'h3a8a3b2b),
	.w6(32'hbae250a9),
	.w7(32'hbb01c59b),
	.w8(32'h3a4fdcb9),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8a6a1b),
	.w1(32'h3a070fef),
	.w2(32'h385a7dec),
	.w3(32'h39b27671),
	.w4(32'h3a1625fe),
	.w5(32'hbacc1c3b),
	.w6(32'h3a33c996),
	.w7(32'h38f3f754),
	.w8(32'hbb9f2c38),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa98b78),
	.w1(32'hbb3bd177),
	.w2(32'hbb30b5d3),
	.w3(32'hbaf49a85),
	.w4(32'hbb02422c),
	.w5(32'h3bf18e53),
	.w6(32'hbc072b44),
	.w7(32'hbb579b88),
	.w8(32'h3c15bc83),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39eed882),
	.w1(32'hbb01fec8),
	.w2(32'h3b0d3447),
	.w3(32'hbb980997),
	.w4(32'h3b3e85e7),
	.w5(32'hbb0323e9),
	.w6(32'hbbb4e2f5),
	.w7(32'h3bc1b623),
	.w8(32'hbb9eb3a1),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab4b62c),
	.w1(32'h3b0f48ad),
	.w2(32'h3b98d103),
	.w3(32'h3b1bbb2a),
	.w4(32'h3b1b87d2),
	.w5(32'hbac40449),
	.w6(32'hbbccfa49),
	.w7(32'h3ab980ee),
	.w8(32'h3a1d467b),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0b276e),
	.w1(32'h37a2f083),
	.w2(32'hbb453712),
	.w3(32'hbb471371),
	.w4(32'h3b5c8f17),
	.w5(32'h3a87f437),
	.w6(32'hbbe67878),
	.w7(32'h3bc2b848),
	.w8(32'h396a071f),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae16ff1),
	.w1(32'hbb13f6a5),
	.w2(32'hbaf51167),
	.w3(32'h3aadcbce),
	.w4(32'hb98b0d7d),
	.w5(32'h3b73603e),
	.w6(32'hba8aad8c),
	.w7(32'h363ab788),
	.w8(32'h3c0ad5a4),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb1341e),
	.w1(32'hb8bb9563),
	.w2(32'h3b9f1480),
	.w3(32'h3b6d7b3a),
	.w4(32'h3bd4b238),
	.w5(32'hba3ce872),
	.w6(32'h3b5c1f43),
	.w7(32'h3bc892a8),
	.w8(32'hbb916267),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0bdb28),
	.w1(32'h3b1c915a),
	.w2(32'hba7a11a1),
	.w3(32'h3ade564c),
	.w4(32'h3b629f3d),
	.w5(32'hba8e13de),
	.w6(32'h39974c1e),
	.w7(32'h3bb3d38d),
	.w8(32'h3b405612),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b82bcb0),
	.w1(32'hba8b9f39),
	.w2(32'hbaf6685b),
	.w3(32'hbc36fe2f),
	.w4(32'hbb7f7343),
	.w5(32'h3c05e703),
	.w6(32'hbaeb90a4),
	.w7(32'hb99e248c),
	.w8(32'h3ab80153),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b860510),
	.w1(32'h3bac0444),
	.w2(32'hbbb66540),
	.w3(32'h3c02505f),
	.w4(32'hbbb7ccfb),
	.w5(32'hbaafcb72),
	.w6(32'hbaff84c9),
	.w7(32'hba259682),
	.w8(32'hbbc2509e),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2c375b),
	.w1(32'h3a3a235c),
	.w2(32'h3bc67a9b),
	.w3(32'hba954f6f),
	.w4(32'h3b8e64e9),
	.w5(32'h3ae2016e),
	.w6(32'hbaeddd8c),
	.w7(32'h3bd47dfa),
	.w8(32'hbaf18dca),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba6f2999),
	.w1(32'hbab1a0c6),
	.w2(32'hbab9054e),
	.w3(32'h3a717fd6),
	.w4(32'h3a1c63ea),
	.w5(32'hbace81b7),
	.w6(32'hbbf14001),
	.w7(32'hbaebbaa3),
	.w8(32'hbb08e174),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0ec736),
	.w1(32'h3b47e89e),
	.w2(32'hbab0488c),
	.w3(32'h39ccf36c),
	.w4(32'hbba849de),
	.w5(32'h3b286dab),
	.w6(32'h3b09cede),
	.w7(32'hbb685466),
	.w8(32'hba6902ed),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9878b5a),
	.w1(32'hbb751cb5),
	.w2(32'hbaf9efc0),
	.w3(32'h3b9af6db),
	.w4(32'h3b2ab4ee),
	.w5(32'h3b9fb205),
	.w6(32'hbacc1c6f),
	.w7(32'h3b7a0b06),
	.w8(32'h3c1d9aa1),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb0a0e7),
	.w1(32'h394e835b),
	.w2(32'hbb0dcad1),
	.w3(32'h3a27cbc3),
	.w4(32'hbb2fcfd7),
	.w5(32'hbb353866),
	.w6(32'h3a32254c),
	.w7(32'hbae1d5a0),
	.w8(32'hbbd3652e),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6d7f5a),
	.w1(32'hbbdaeff1),
	.w2(32'hbbf1ed04),
	.w3(32'hbb7c7da0),
	.w4(32'hbba46d2b),
	.w5(32'hba24cd0b),
	.w6(32'hbbad4ce3),
	.w7(32'hbc13bfa5),
	.w8(32'hba6f13fa),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3490f9),
	.w1(32'hba4f935b),
	.w2(32'hb9b9d220),
	.w3(32'h39e03b7a),
	.w4(32'hbb5fe0e7),
	.w5(32'hbbcfc19c),
	.w6(32'hbb462196),
	.w7(32'hbba754cb),
	.w8(32'hbbf4597d),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb94cd76),
	.w1(32'hbbdd7b8f),
	.w2(32'h3ae0ae42),
	.w3(32'hbbb76260),
	.w4(32'hba6a2ed9),
	.w5(32'hbb70a6de),
	.w6(32'hbb970027),
	.w7(32'h39860c82),
	.w8(32'hb9fe13dd),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3af12b37),
	.w1(32'h3a8961b8),
	.w2(32'h3a157094),
	.w3(32'h3ae66025),
	.w4(32'hbad9e437),
	.w5(32'hbac43eb6),
	.w6(32'h39640f54),
	.w7(32'h39b5c39f),
	.w8(32'hba8c490b),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadbaa6b),
	.w1(32'hbaa5de56),
	.w2(32'hbb9021c9),
	.w3(32'hbaad2280),
	.w4(32'hbb7fbe08),
	.w5(32'h39cb3768),
	.w6(32'hbadc76a8),
	.w7(32'hbb865f02),
	.w8(32'h3b471f38),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4ece85),
	.w1(32'h3b19007b),
	.w2(32'hbb990286),
	.w3(32'hbb95ada7),
	.w4(32'h3b430404),
	.w5(32'h3b28dc84),
	.w6(32'hb6ae297f),
	.w7(32'h3ac33d2c),
	.w8(32'h3a517957),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac9e9aa),
	.w1(32'hba85e1f5),
	.w2(32'h3b1aedcb),
	.w3(32'h3b10d7bc),
	.w4(32'h3b06653b),
	.w5(32'hbbc5ed51),
	.w6(32'hbad1712f),
	.w7(32'h3b5cd5ee),
	.w8(32'hbc4cf529),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc463101),
	.w1(32'hbc536426),
	.w2(32'hbbadb89c),
	.w3(32'hbba0c41c),
	.w4(32'hbb4ccdf1),
	.w5(32'h3b0d7601),
	.w6(32'hbc6c3c8f),
	.w7(32'hbba2cd4c),
	.w8(32'h3ae671b4),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b047485),
	.w1(32'h399e0dbd),
	.w2(32'h3b7b46d2),
	.w3(32'h3c0200af),
	.w4(32'hba966035),
	.w5(32'h3ad54e1b),
	.w6(32'h3bf1dde9),
	.w7(32'hbb07bd30),
	.w8(32'hbb43c13d),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb894dc73),
	.w1(32'h3bb7b856),
	.w2(32'hbbd25930),
	.w3(32'h3b920364),
	.w4(32'hbb6875c0),
	.w5(32'h3b43b840),
	.w6(32'h3c277ed9),
	.w7(32'hbb974ff0),
	.w8(32'h3a483e3e),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2fe288),
	.w1(32'hbbb3742a),
	.w2(32'hbb764de0),
	.w3(32'h3aa65201),
	.w4(32'h3b6bb728),
	.w5(32'h3bab3092),
	.w6(32'hbbfcbf31),
	.w7(32'hbb5eb9f6),
	.w8(32'h3b18e902),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9dc0fa),
	.w1(32'h39161587),
	.w2(32'hbbb61e36),
	.w3(32'hbb91bb77),
	.w4(32'hbb56ca86),
	.w5(32'h3ba4103b),
	.w6(32'h3b6e9ae9),
	.w7(32'hbbcfca36),
	.w8(32'h3b3ed2f8),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b687283),
	.w1(32'hbb6f3deb),
	.w2(32'h3b27f0e1),
	.w3(32'h3b2c9f22),
	.w4(32'hbaf04fe8),
	.w5(32'hba01b52d),
	.w6(32'h3ae39135),
	.w7(32'hbaedb727),
	.w8(32'h3b68c2ef),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b009fa5),
	.w1(32'h3aaf6c10),
	.w2(32'hbba7225e),
	.w3(32'hbadd1581),
	.w4(32'h3b85db68),
	.w5(32'h38ce2860),
	.w6(32'h3ae61997),
	.w7(32'hba664d4e),
	.w8(32'hbad55f0e),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb236b37),
	.w1(32'h3b22106e),
	.w2(32'h3b92b6b9),
	.w3(32'h3a766dad),
	.w4(32'hba4726d1),
	.w5(32'h3ae7c2e8),
	.w6(32'h3af8a0b2),
	.w7(32'h3b05cffe),
	.w8(32'h3acd6b8f),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39087d8e),
	.w1(32'hb9752818),
	.w2(32'hbb04c7c7),
	.w3(32'h3b64ed6e),
	.w4(32'hba7c3574),
	.w5(32'hbba81974),
	.w6(32'h3b33d9f4),
	.w7(32'hbb73fa03),
	.w8(32'hbacfecf0),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2d3a85),
	.w1(32'h3b4cae4b),
	.w2(32'hbb0aa535),
	.w3(32'hb90716b3),
	.w4(32'hbb4aa2b8),
	.w5(32'h3ad6d651),
	.w6(32'h3b74a493),
	.w7(32'hbb30a507),
	.w8(32'hbbf439fa),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb236c0b),
	.w1(32'hbad2867f),
	.w2(32'h3a803963),
	.w3(32'hbb42b418),
	.w4(32'h3947abe3),
	.w5(32'hbb9c9135),
	.w6(32'hbb49d8f3),
	.w7(32'hbb248f9d),
	.w8(32'hbbb87f49),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7f1547),
	.w1(32'h3b3c61d3),
	.w2(32'hba7f51af),
	.w3(32'h3c1b0410),
	.w4(32'h3b54657b),
	.w5(32'hba626076),
	.w6(32'h3b9e491e),
	.w7(32'h39e23b56),
	.w8(32'hbb128866),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4a8831),
	.w1(32'hbab50080),
	.w2(32'hbac91323),
	.w3(32'h3a728e10),
	.w4(32'h3a659dd7),
	.w5(32'hbbb700c5),
	.w6(32'hbb562608),
	.w7(32'h3b52cc34),
	.w8(32'h3a9519cc),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc682d8),
	.w1(32'hbbe43b76),
	.w2(32'hbbdeafe9),
	.w3(32'hbba44cae),
	.w4(32'hbbe08fe1),
	.w5(32'hbae7cddb),
	.w6(32'hbb933967),
	.w7(32'h3b84c8c4),
	.w8(32'hbb750644),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb21b726),
	.w1(32'hba42a7ba),
	.w2(32'hba1ed25a),
	.w3(32'hba25b73d),
	.w4(32'hbabb5f28),
	.w5(32'h3a6cf8f9),
	.w6(32'hbae0b7fb),
	.w7(32'hbac23553),
	.w8(32'hbb17b8d7),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a934cd),
	.w1(32'hb99d415f),
	.w2(32'hbab7cca2),
	.w3(32'h384e44ac),
	.w4(32'hbb0904e0),
	.w5(32'hbbce6ba5),
	.w6(32'hbafa698e),
	.w7(32'hbacd297e),
	.w8(32'hbb40a2ef),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb47ef5c),
	.w1(32'hbbb3fafd),
	.w2(32'hbc359105),
	.w3(32'hbbf6e970),
	.w4(32'hbb9a6335),
	.w5(32'hbb4ce869),
	.w6(32'hbc02eb05),
	.w7(32'hbbb1151a),
	.w8(32'hbb95fe8c),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4e51a8),
	.w1(32'hbb624529),
	.w2(32'hbbb1d4c8),
	.w3(32'hbba24958),
	.w4(32'hbbc601c4),
	.w5(32'hb9ac87ad),
	.w6(32'hbb919b62),
	.w7(32'hbbbd3782),
	.w8(32'hbb016b81),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaa7221),
	.w1(32'hb9bc6528),
	.w2(32'h391375ce),
	.w3(32'h3a0c2834),
	.w4(32'hba579518),
	.w5(32'hbbbe4448),
	.w6(32'hba8faaae),
	.w7(32'hb9b1f599),
	.w8(32'hbbced8d8),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb80bc13),
	.w1(32'hbb0c90aa),
	.w2(32'h3ae7be56),
	.w3(32'h37757700),
	.w4(32'h3b9c1509),
	.w5(32'h3bad9765),
	.w6(32'hbb514a79),
	.w7(32'h3b35472d),
	.w8(32'hbaec40c9),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b88c0f3),
	.w1(32'h3b833110),
	.w2(32'hb9089dd2),
	.w3(32'h3bcc53e6),
	.w4(32'hbab3f798),
	.w5(32'h3bbf7d90),
	.w6(32'h3a661193),
	.w7(32'hbb2a6883),
	.w8(32'h3c21b561),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba65ca8),
	.w1(32'hbbaac9a1),
	.w2(32'hbc420d2e),
	.w3(32'hbbac85f2),
	.w4(32'hbc13f5cf),
	.w5(32'hbaaf85c3),
	.w6(32'hbb0bc352),
	.w7(32'hbbd1de1b),
	.w8(32'h3c04fe1f),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b570d86),
	.w1(32'h3a82cedf),
	.w2(32'hba69703c),
	.w3(32'hbb901c69),
	.w4(32'h37eac602),
	.w5(32'h3a962e32),
	.w6(32'h3a09f21e),
	.w7(32'h3ac8510c),
	.w8(32'hba0167d0),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b02af0c),
	.w1(32'hba8004c5),
	.w2(32'hba25bc5e),
	.w3(32'h3b4b708b),
	.w4(32'h3b7a95cf),
	.w5(32'h3b136c51),
	.w6(32'h39d27727),
	.w7(32'h3b4a0edd),
	.w8(32'hbaa59e65),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae356e2),
	.w1(32'hbb1f889e),
	.w2(32'h3b6d9639),
	.w3(32'hb8cd3fe2),
	.w4(32'h3bfbed3a),
	.w5(32'h3b0109ee),
	.w6(32'hbb1b37bf),
	.w7(32'h3bf29063),
	.w8(32'hba370e86),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39cbedf9),
	.w1(32'hbafbaab0),
	.w2(32'h3a310c9a),
	.w3(32'hbb0aeacd),
	.w4(32'hba309993),
	.w5(32'h394dc39c),
	.w6(32'hbb19c368),
	.w7(32'hba499cd7),
	.w8(32'h3b487659),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b327370),
	.w1(32'hbb316a61),
	.w2(32'hbb710c73),
	.w3(32'hbb5e2414),
	.w4(32'hbb8e7c95),
	.w5(32'hba016690),
	.w6(32'h39b37f83),
	.w7(32'hbb7e7ec9),
	.w8(32'h3b82ea8b),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb708d5a),
	.w1(32'hbbcb83f2),
	.w2(32'h3b8ca9dc),
	.w3(32'hbad77bce),
	.w4(32'h3b23cf19),
	.w5(32'h3bc057a3),
	.w6(32'hbae17388),
	.w7(32'h3b5345fc),
	.w8(32'h3acbe867),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb32b8ba),
	.w1(32'h3ae9db3c),
	.w2(32'hbad9bf4f),
	.w3(32'hbb6510fd),
	.w4(32'hbbc2b159),
	.w5(32'hbb81b89a),
	.w6(32'h3bf50d35),
	.w7(32'hbbbb7f13),
	.w8(32'hbbe62239),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb943a0b),
	.w1(32'hbb05a206),
	.w2(32'h3bc5c119),
	.w3(32'hbb99de97),
	.w4(32'h3c463a15),
	.w5(32'hbb05624b),
	.w6(32'hbb821154),
	.w7(32'h3c1181b4),
	.w8(32'hbb69ce6a),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb656b28),
	.w1(32'hbb90f792),
	.w2(32'hbb4648a4),
	.w3(32'h3a819104),
	.w4(32'hb9f1f7da),
	.w5(32'h3ae01ff0),
	.w6(32'hbb70dd12),
	.w7(32'hba8231c4),
	.w8(32'hba9ae6d0),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb990722a),
	.w1(32'hbb192fd7),
	.w2(32'hb9ee093d),
	.w3(32'h3b8d5cb2),
	.w4(32'hb97b1612),
	.w5(32'h3998021e),
	.w6(32'h3af93116),
	.w7(32'hbac9b91d),
	.w8(32'hbb89a2b2),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb87b156),
	.w1(32'h3afadf47),
	.w2(32'h3aa8c1a2),
	.w3(32'h3b8709eb),
	.w4(32'h3bf957aa),
	.w5(32'hbbaf42dd),
	.w6(32'h3ae4c7ad),
	.w7(32'h3c52ef92),
	.w8(32'hbb3e116a),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba85cb12),
	.w1(32'hbaf71676),
	.w2(32'hbb8f298b),
	.w3(32'hbae8a6e9),
	.w4(32'hbb2c1ee9),
	.w5(32'h3ada9d55),
	.w6(32'hbbae3f6b),
	.w7(32'hbb155131),
	.w8(32'h3b2811b8),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b7ad5c2),
	.w1(32'hba868608),
	.w2(32'h3b2e4462),
	.w3(32'h3b02c106),
	.w4(32'h3b4d8c28),
	.w5(32'h3b43ebdd),
	.w6(32'hba65fd85),
	.w7(32'h3b4818b0),
	.w8(32'hba4af7ba),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0c8c18),
	.w1(32'h3a08be61),
	.w2(32'hb9a50d05),
	.w3(32'h3ba923d5),
	.w4(32'h3b361a41),
	.w5(32'hba6f4c4b),
	.w6(32'hbae57dbc),
	.w7(32'hb8799f5d),
	.w8(32'hbb0050b9),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5464eb),
	.w1(32'h36ae8956),
	.w2(32'hbb028140),
	.w3(32'hbaf684b4),
	.w4(32'hbbc27b5c),
	.w5(32'h3b31910e),
	.w6(32'h38b42a1b),
	.w7(32'hbb7e314b),
	.w8(32'h3bdd0411),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8e80f8),
	.w1(32'h3bb5ef0e),
	.w2(32'hbbe3a035),
	.w3(32'hbc025943),
	.w4(32'h3b6d3b9d),
	.w5(32'h3c159125),
	.w6(32'hbb1de23f),
	.w7(32'hbaa0c43f),
	.w8(32'h3bb87135),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b485da2),
	.w1(32'h3bd7b162),
	.w2(32'hbb0c657a),
	.w3(32'h3c210236),
	.w4(32'hbb275128),
	.w5(32'hb9e5fa8b),
	.w6(32'h3c70c9ce),
	.w7(32'hbb33da99),
	.w8(32'hbb0c9533),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb58a67a),
	.w1(32'hbb0c1b87),
	.w2(32'hbb421ab3),
	.w3(32'hbbfa6977),
	.w4(32'h3b01829e),
	.w5(32'hbb62f3a9),
	.w6(32'hbb6cbe5e),
	.w7(32'h3c2cebe7),
	.w8(32'hbb19fa3a),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7bab70),
	.w1(32'hbb420d3b),
	.w2(32'hbb24861d),
	.w3(32'hbbcea1f5),
	.w4(32'hb92f28e9),
	.w5(32'h3b694d3b),
	.w6(32'hbafec849),
	.w7(32'h3af0bdb0),
	.w8(32'h3c036603),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba56fb53),
	.w1(32'hbbc30aa6),
	.w2(32'hba36155f),
	.w3(32'h3b2fec3a),
	.w4(32'h3b4398af),
	.w5(32'h3ab66133),
	.w6(32'hbaa55b73),
	.w7(32'h3b86069d),
	.w8(32'h3b2edf34),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b26e831),
	.w1(32'h3bb7074c),
	.w2(32'hbbcf60a5),
	.w3(32'h38c2c807),
	.w4(32'hbbe1b47d),
	.w5(32'hba9f6754),
	.w6(32'h3bb56084),
	.w7(32'hbbd733ca),
	.w8(32'h3abf8b6a),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbafcc6d8),
	.w1(32'h3a194b63),
	.w2(32'hbb970c9a),
	.w3(32'hbb04faa6),
	.w4(32'hba2562f1),
	.w5(32'h3ba5b494),
	.w6(32'h3b9b94cd),
	.w7(32'hbb474b8c),
	.w8(32'hba6b6c53),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac03a2e),
	.w1(32'hbb2137a1),
	.w2(32'h3b98d972),
	.w3(32'hbc13b194),
	.w4(32'h3b25b489),
	.w5(32'hbad60a77),
	.w6(32'hbba6228f),
	.w7(32'h3bb8c972),
	.w8(32'h3b4f4f29),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab776dc),
	.w1(32'hbae7bfb5),
	.w2(32'hbaace9b2),
	.w3(32'hbb3fb1f4),
	.w4(32'h3b96731b),
	.w5(32'hba895e59),
	.w6(32'h3be8e1cb),
	.w7(32'h3b39ded1),
	.w8(32'hba5262e7),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8cc536),
	.w1(32'hbb701835),
	.w2(32'h391c0768),
	.w3(32'h3b6ad534),
	.w4(32'h3acfa73d),
	.w5(32'h3acd321c),
	.w6(32'hbb446d09),
	.w7(32'h3a91dc7e),
	.w8(32'h3b47c95d),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba277a6),
	.w1(32'h3a080439),
	.w2(32'hb9445fb9),
	.w3(32'hbb4e8a5a),
	.w4(32'hbb5871a2),
	.w5(32'hbab8577f),
	.w6(32'h3b78fd34),
	.w7(32'hba4c8b65),
	.w8(32'hbadaddff),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaed9767),
	.w1(32'h3ba9d7c6),
	.w2(32'h3bba3750),
	.w3(32'h3bbc29c8),
	.w4(32'h3b87b25f),
	.w5(32'h3b94f9e2),
	.w6(32'h3bf27306),
	.w7(32'h3ba0fe89),
	.w8(32'h3be211d5),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b94b2bd),
	.w1(32'h3c09bb3b),
	.w2(32'hbb40cc81),
	.w3(32'hba38533c),
	.w4(32'hbb97eb12),
	.w5(32'h394979fd),
	.w6(32'h3bd62d22),
	.w7(32'hbbc23d68),
	.w8(32'h39b2eaf7),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a1ef7ce),
	.w1(32'h3a8a1b70),
	.w2(32'h3b7c038e),
	.w3(32'h3b3c951e),
	.w4(32'h3a641edc),
	.w5(32'hbbec1429),
	.w6(32'hba111457),
	.w7(32'h3b48a622),
	.w8(32'hbbb24e5d),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb853e16),
	.w1(32'hbb30d839),
	.w2(32'h3b4da9c9),
	.w3(32'hba49787c),
	.w4(32'h3a8c5182),
	.w5(32'h3bb4b7a0),
	.w6(32'hb9095844),
	.w7(32'hb9b6c713),
	.w8(32'hbbeae1dd),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39da9900),
	.w1(32'h3aa56123),
	.w2(32'h3c1b3f48),
	.w3(32'h3ac0773f),
	.w4(32'h3c3aeb37),
	.w5(32'hbc1ab250),
	.w6(32'hbb95251c),
	.w7(32'h3c3a4658),
	.w8(32'hbc1226f8),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc005706),
	.w1(32'hbc569ccf),
	.w2(32'hba930ea0),
	.w3(32'hbba20133),
	.w4(32'hba8a336f),
	.w5(32'h3a3b2e6f),
	.w6(32'hbc81c367),
	.w7(32'hb9f1b5b8),
	.w8(32'hb99f3898),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2289ae),
	.w1(32'h3c29f028),
	.w2(32'hba9282fa),
	.w3(32'h3afd7c64),
	.w4(32'hbbd07fb9),
	.w5(32'hba641981),
	.w6(32'h3ba02217),
	.w7(32'hbb35854b),
	.w8(32'hbbdbe1e8),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb93b08ad),
	.w1(32'h3b4f009a),
	.w2(32'hbb40955d),
	.w3(32'h3a7a58a9),
	.w4(32'hbadf41e1),
	.w5(32'hbabc43ad),
	.w6(32'hbb742c11),
	.w7(32'hbb5b9387),
	.w8(32'hbb7e32ba),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6a0b83),
	.w1(32'hbbf3d2a6),
	.w2(32'hbbfe4677),
	.w3(32'hbb05ceb7),
	.w4(32'hbb13e7dc),
	.w5(32'h3a46f961),
	.w6(32'hbb9c3180),
	.w7(32'hbb9ae7e1),
	.w8(32'h3919ddcb),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38dfaa5f),
	.w1(32'hbb562bfa),
	.w2(32'hbbc2630b),
	.w3(32'hbbbe5619),
	.w4(32'hbbc2ca68),
	.w5(32'h3a8a9c2c),
	.w6(32'hbb0382bd),
	.w7(32'hbb71efed),
	.w8(32'hbab49359),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1d1624),
	.w1(32'hbb7a3d9a),
	.w2(32'hbb1808b8),
	.w3(32'h3b9f485f),
	.w4(32'h3a9ce68e),
	.w5(32'h3ab440ce),
	.w6(32'hba5f70b8),
	.w7(32'h39dc4797),
	.w8(32'h3b066e31),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad26e7d),
	.w1(32'hb915dcc8),
	.w2(32'hbab0a5a0),
	.w3(32'h3b2f2a86),
	.w4(32'hbb49fa43),
	.w5(32'h3a438824),
	.w6(32'hba042b58),
	.w7(32'h391e373f),
	.w8(32'h3a3c31dd),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9188ef),
	.w1(32'hbb2f2c35),
	.w2(32'h3a7c7e6f),
	.w3(32'hbba291e7),
	.w4(32'h3b6329d8),
	.w5(32'hbaa874cb),
	.w6(32'hbb384372),
	.w7(32'h3ae487fc),
	.w8(32'h39a6dd8c),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae551f2),
	.w1(32'hbaa9bb9a),
	.w2(32'h3b7b0cc6),
	.w3(32'h3b974775),
	.w4(32'hba03c958),
	.w5(32'h3b890804),
	.w6(32'h3aac1d20),
	.w7(32'h3af13a0d),
	.w8(32'hbacb23a5),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa3fed7),
	.w1(32'h3c500071),
	.w2(32'hbc221c59),
	.w3(32'h3ca29cd3),
	.w4(32'hbc0f28c9),
	.w5(32'h3b36bd7d),
	.w6(32'h3cc8e217),
	.w7(32'hbc9b1d44),
	.w8(32'hba6e5c6b),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb363781),
	.w1(32'h3a23cdf5),
	.w2(32'h3b71afdb),
	.w3(32'hba983ce0),
	.w4(32'h3a83e31d),
	.w5(32'hbb7beed7),
	.w6(32'h3b6973dc),
	.w7(32'hb90e63fa),
	.w8(32'hbb1f575c),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb74c433),
	.w1(32'hbb1b8e8d),
	.w2(32'hb9fee04f),
	.w3(32'hbbbdae0f),
	.w4(32'h3ad3d1fd),
	.w5(32'hbb533de6),
	.w6(32'hbb95ae0e),
	.w7(32'h3b8da512),
	.w8(32'h3abab744),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba75dbaf),
	.w1(32'h3a882204),
	.w2(32'hbb40b843),
	.w3(32'hbc05cc17),
	.w4(32'hbb33edf9),
	.w5(32'hba5b60a9),
	.w6(32'hb9a2b7e3),
	.w7(32'hbb720a10),
	.w8(32'hbb24b7b0),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2bf544),
	.w1(32'h3b07fc78),
	.w2(32'hba8823f7),
	.w3(32'hb9843fc2),
	.w4(32'hbae0c466),
	.w5(32'hb9be37da),
	.w6(32'h3ae81530),
	.w7(32'hbb2a1f86),
	.w8(32'hbaa5ee40),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb472a28),
	.w1(32'hbb0a5bbc),
	.w2(32'hbb4a0592),
	.w3(32'h3b67384d),
	.w4(32'h385f660d),
	.w5(32'hbc23a89a),
	.w6(32'hbaea2adb),
	.w7(32'hbaa275e3),
	.w8(32'hbc06fb04),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2e2e2b),
	.w1(32'hbc6b329f),
	.w2(32'hbbe02b07),
	.w3(32'hbc268400),
	.w4(32'hbbb10ed4),
	.w5(32'hb9e1c37b),
	.w6(32'hbc54f085),
	.w7(32'hbb86bc41),
	.w8(32'hb9193e22),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3ddb4d),
	.w1(32'h392aafac),
	.w2(32'h39d8461a),
	.w3(32'h3ae0fb81),
	.w4(32'hba1eeeb2),
	.w5(32'h3ae59d86),
	.w6(32'h3b797514),
	.w7(32'h3ae8abaa),
	.w8(32'h3aaa116c),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7ce988),
	.w1(32'h3b479b69),
	.w2(32'h3b784b29),
	.w3(32'h3b957a8a),
	.w4(32'h393d5d01),
	.w5(32'hbb4904f7),
	.w6(32'h3b827177),
	.w7(32'h3b82017c),
	.w8(32'hba7d0006),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb695eb7),
	.w1(32'hbb08dbf3),
	.w2(32'h3b603ef1),
	.w3(32'hbb963fcb),
	.w4(32'hbbb20d0e),
	.w5(32'h3b962d9f),
	.w6(32'hbad69a38),
	.w7(32'hbb5412f0),
	.w8(32'h3bf11d43),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb3a5d4),
	.w1(32'h3c03be39),
	.w2(32'hbb53049b),
	.w3(32'hbad7b512),
	.w4(32'h38325f1b),
	.w5(32'h3c17f451),
	.w6(32'h3c0ccf8e),
	.w7(32'hba75e5a0),
	.w8(32'h3c076f25),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9ccf82),
	.w1(32'h3bf53b17),
	.w2(32'h3a48408b),
	.w3(32'h3c0af840),
	.w4(32'hba1a8b9c),
	.w5(32'hbb858fbc),
	.w6(32'h3c93f911),
	.w7(32'hb97e2af5),
	.w8(32'hbbaaef25),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb90e0bf),
	.w1(32'hbbc6c3c7),
	.w2(32'h3b6438a5),
	.w3(32'h3b5a439b),
	.w4(32'h39b7d25a),
	.w5(32'hbbb2fe13),
	.w6(32'hbb74377e),
	.w7(32'hba7bb377),
	.w8(32'hbaa4153c),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7ab2f8),
	.w1(32'h3ac9302b),
	.w2(32'hbbb6b0cd),
	.w3(32'hbad70c7e),
	.w4(32'h38dba564),
	.w5(32'h39a59f42),
	.w6(32'h3a742e30),
	.w7(32'hbb486141),
	.w8(32'hbb79efdf),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1a5842),
	.w1(32'hbb93bd7e),
	.w2(32'hbae22148),
	.w3(32'hbb8690e9),
	.w4(32'h3a98dfe5),
	.w5(32'hbb8facc0),
	.w6(32'hbbb34d31),
	.w7(32'h3ac44db6),
	.w8(32'hbbc93721),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcd04fd),
	.w1(32'h3b014d8b),
	.w2(32'hba9dc85f),
	.w3(32'h3ab1a6c6),
	.w4(32'hbb0b6152),
	.w5(32'h3b022c42),
	.w6(32'h3b369aa8),
	.w7(32'hbb331e71),
	.w8(32'hba3ee0c5),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8a8fe7),
	.w1(32'h3b97c54f),
	.w2(32'hbb3a01d3),
	.w3(32'hbb7ca32f),
	.w4(32'hbb3fce58),
	.w5(32'hbba8d65d),
	.w6(32'h39708067),
	.w7(32'h396ed7fc),
	.w8(32'hbbb4fade),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb35b919),
	.w1(32'hbbb639d9),
	.w2(32'h3b604519),
	.w3(32'hbad0c5c6),
	.w4(32'h3b70176a),
	.w5(32'h3bb053cb),
	.w6(32'hbbc68f1f),
	.w7(32'h3b941e42),
	.w8(32'hbaa6d806),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbabaf3ce),
	.w1(32'h3b3c4c1c),
	.w2(32'h3bc6ac6d),
	.w3(32'hbb7b50fb),
	.w4(32'h3b819cfc),
	.w5(32'hba8fdcdc),
	.w6(32'hbb45f116),
	.w7(32'h3c3413cc),
	.w8(32'h3b43434c),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h385a125d),
	.w1(32'hbaa6bb3e),
	.w2(32'hbaae2ca8),
	.w3(32'hbb004ef8),
	.w4(32'hba2d82f7),
	.w5(32'h3c29ab85),
	.w6(32'hbb591212),
	.w7(32'h3b60b809),
	.w8(32'h3c247cea),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baeb087),
	.w1(32'h3bd49783),
	.w2(32'hbb71330d),
	.w3(32'hbb7f121d),
	.w4(32'hbbcf707c),
	.w5(32'hbb5d3dff),
	.w6(32'h3c54f05d),
	.w7(32'hbbd01f15),
	.w8(32'hbb88a3c6),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1dd6db),
	.w1(32'h3a9a490b),
	.w2(32'hba2b9499),
	.w3(32'h3b101226),
	.w4(32'h3b1e96ff),
	.w5(32'h3afc5c8b),
	.w6(32'h3bb8512c),
	.w7(32'hbb051117),
	.w8(32'h3bcc96de),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b429e87),
	.w1(32'hba531222),
	.w2(32'hbb98ef56),
	.w3(32'hbc152f1c),
	.w4(32'hbbaf1fc9),
	.w5(32'hba80b06a),
	.w6(32'hba986bd2),
	.w7(32'hbb68e4e1),
	.w8(32'hbb390209),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1aee85),
	.w1(32'hbbacdbf0),
	.w2(32'h3b33efd0),
	.w3(32'h3aa2c832),
	.w4(32'hba108ef9),
	.w5(32'hb803dc1d),
	.w6(32'hbbf58c0d),
	.w7(32'hba08b3a9),
	.w8(32'hba98844d),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc3f710),
	.w1(32'hba9f3453),
	.w2(32'h364bdd2c),
	.w3(32'hbb29b7f7),
	.w4(32'h3b000bd9),
	.w5(32'h3b99fb13),
	.w6(32'hbc137c0a),
	.w7(32'hb9e83b34),
	.w8(32'h3c057969),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3f27c1),
	.w1(32'hb9232f9f),
	.w2(32'hbb1d0479),
	.w3(32'hbb1aad6b),
	.w4(32'h39fe7fa2),
	.w5(32'hbaa4c216),
	.w6(32'h391b3c86),
	.w7(32'h3b05e2de),
	.w8(32'hbb8cbfae),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4511ea),
	.w1(32'hbab5c22a),
	.w2(32'hbb6ff664),
	.w3(32'hbb881ec4),
	.w4(32'hbb8dd138),
	.w5(32'hbc01c076),
	.w6(32'hbb5a74ea),
	.w7(32'hbbbe9fdb),
	.w8(32'hbbb30f56),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc04e1f3),
	.w1(32'hbb090134),
	.w2(32'hbae4e969),
	.w3(32'hbbefbe86),
	.w4(32'h3a660766),
	.w5(32'hba709c23),
	.w6(32'hbb37f544),
	.w7(32'h3bb4caa3),
	.w8(32'h3bd36aa9),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b718cb3),
	.w1(32'hba2106c9),
	.w2(32'hbb4da77e),
	.w3(32'hbba55442),
	.w4(32'hbbdc2db7),
	.w5(32'hbb55fc79),
	.w6(32'h3b958d65),
	.w7(32'hbb4d8a5f),
	.w8(32'hbb3e30df),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f98539),
	.w1(32'h3b8fdc5b),
	.w2(32'h3a927724),
	.w3(32'h3be3453e),
	.w4(32'h3a8791ec),
	.w5(32'h3bbc11e0),
	.w6(32'h3c29e863),
	.w7(32'h3bcaa514),
	.w8(32'h3aed7b44),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b11643d),
	.w1(32'h3bba8f38),
	.w2(32'h3bb54b88),
	.w3(32'h3bbf121d),
	.w4(32'h3bfde0be),
	.w5(32'hbb4eb36a),
	.w6(32'h3af00109),
	.w7(32'h3c4246be),
	.w8(32'hbbc63d2b),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb76251b6),
	.w1(32'h3b69df8b),
	.w2(32'h3a183369),
	.w3(32'h3b945242),
	.w4(32'h393eb2b4),
	.w5(32'hbb4a347c),
	.w6(32'h3b97cbe4),
	.w7(32'h3b5c9fd3),
	.w8(32'hba181fac),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb465051),
	.w1(32'h3aea8b2c),
	.w2(32'h3b156b2f),
	.w3(32'h3ad52b22),
	.w4(32'h3a88beff),
	.w5(32'h3b6111b6),
	.w6(32'hba6a3029),
	.w7(32'h3b89b004),
	.w8(32'hbc00e564),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a684706),
	.w1(32'h3bd240e8),
	.w2(32'hba9f0713),
	.w3(32'h3c12a01e),
	.w4(32'h3baaa9a3),
	.w5(32'hba9c5a98),
	.w6(32'h3b3393b6),
	.w7(32'h3a493002),
	.w8(32'hbb796410),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc70496),
	.w1(32'hbb8c75a9),
	.w2(32'hbb23a513),
	.w3(32'hba9f9c10),
	.w4(32'h38ea78c3),
	.w5(32'h3a0722d8),
	.w6(32'hbaaa8b55),
	.w7(32'hbab629f2),
	.w8(32'hbb1dd2ed),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9a6caa),
	.w1(32'hbb370f82),
	.w2(32'hbb10dae5),
	.w3(32'hb9e156b3),
	.w4(32'hbb34343e),
	.w5(32'h38de81e5),
	.w6(32'hbad57370),
	.w7(32'hbb0066e1),
	.w8(32'h3a485f1f),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab85f61),
	.w1(32'h3899c507),
	.w2(32'hbc0eff3d),
	.w3(32'hbbc5b18c),
	.w4(32'hbb9c8439),
	.w5(32'hbaaf33ac),
	.w6(32'hbb0f1aee),
	.w7(32'hbc1bb398),
	.w8(32'hbbbf8bd1),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb00e9f5),
	.w1(32'h3be11ee3),
	.w2(32'h3b568dab),
	.w3(32'h3c37e59d),
	.w4(32'hbb3e2d69),
	.w5(32'h3b4ed294),
	.w6(32'h3c0bbb15),
	.w7(32'h3a658306),
	.w8(32'h3bfd3e1d),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a3cd92a),
	.w1(32'hbb0a15e8),
	.w2(32'hbb131a45),
	.w3(32'hba4e448c),
	.w4(32'hbb4c16ae),
	.w5(32'hbb56c6ab),
	.w6(32'hbb068314),
	.w7(32'hbb0a1563),
	.w8(32'hbb97c601),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb6cf25),
	.w1(32'hbb38c9b9),
	.w2(32'h3bdc498e),
	.w3(32'h3a2da184),
	.w4(32'h3b9667e8),
	.w5(32'h3b925733),
	.w6(32'hbb36bf01),
	.w7(32'h3a8b3d6d),
	.w8(32'h3a4bf08e),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae0a679),
	.w1(32'h3b2a9122),
	.w2(32'hbaee835e),
	.w3(32'h3b9e6783),
	.w4(32'hb9ee7494),
	.w5(32'h39ce4074),
	.w6(32'h3b075164),
	.w7(32'hbae6a62a),
	.w8(32'h3a2e9c70),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aef5593),
	.w1(32'hbaff46c3),
	.w2(32'h3c00fdb3),
	.w3(32'h3a0f2a93),
	.w4(32'h3bb532a3),
	.w5(32'hbb0dbc09),
	.w6(32'hbb4c1e83),
	.w7(32'h3bf237e8),
	.w8(32'hbb679365),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9e22d4),
	.w1(32'hbba6924e),
	.w2(32'h3af18214),
	.w3(32'hba21ba0e),
	.w4(32'h3bdfef2a),
	.w5(32'h3bbcccb9),
	.w6(32'hbbfc5cb3),
	.w7(32'h3b694454),
	.w8(32'h3c204f45),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba96d58),
	.w1(32'hb83108fe),
	.w2(32'h3ba2e98b),
	.w3(32'hb956d8db),
	.w4(32'h3ac1dba5),
	.w5(32'hb7a53cb7),
	.w6(32'h3b517ffa),
	.w7(32'h3bb0617d),
	.w8(32'hba84d13b),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0532ad),
	.w1(32'hbc1697a5),
	.w2(32'hb90fd595),
	.w3(32'hbbb29e0a),
	.w4(32'hbaf138f1),
	.w5(32'hb9640d0d),
	.w6(32'hbb99f5dc),
	.w7(32'h3b583bee),
	.w8(32'hb9633432),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398b8f88),
	.w1(32'hba52e0ea),
	.w2(32'hb9b14943),
	.w3(32'hb932cab4),
	.w4(32'hb9608921),
	.w5(32'hbb1626d0),
	.w6(32'hba8bb66c),
	.w7(32'hba110731),
	.w8(32'hbb193d64),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b18e837),
	.w1(32'hba75b3ef),
	.w2(32'hba2250fa),
	.w3(32'hbb36345a),
	.w4(32'hb9c5984a),
	.w5(32'h39394026),
	.w6(32'hbaab85c5),
	.w7(32'hba99ead0),
	.w8(32'hba589bb1),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a27f95c),
	.w1(32'hb85134f2),
	.w2(32'hba98a329),
	.w3(32'hbac44926),
	.w4(32'hbac9e1ea),
	.w5(32'h3aaaed08),
	.w6(32'hbb267b22),
	.w7(32'hbb3162fc),
	.w8(32'h3aa04693),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39eaf3b9),
	.w1(32'h3aaa662c),
	.w2(32'h3b181061),
	.w3(32'hbaa37b83),
	.w4(32'hbb103991),
	.w5(32'hbb0df58c),
	.w6(32'h3a7ea70b),
	.w7(32'h39cb6cf9),
	.w8(32'hbabaa6a4),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ca8d9c),
	.w1(32'h3b863085),
	.w2(32'h39cb63af),
	.w3(32'h39e14f10),
	.w4(32'h3b3629b2),
	.w5(32'hbb4caf31),
	.w6(32'h3b837e0d),
	.w7(32'h3b10710b),
	.w8(32'hbb565aed),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba14304b),
	.w1(32'hbab00e98),
	.w2(32'hbb6cfed8),
	.w3(32'hbb0aac19),
	.w4(32'hbb889b57),
	.w5(32'h3abf9d77),
	.w6(32'hbb2c40ae),
	.w7(32'hbb71d8d5),
	.w8(32'h3b0933a3),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38ac5bcf),
	.w1(32'hb904b1a8),
	.w2(32'hbb347d33),
	.w3(32'hba98cb63),
	.w4(32'hba17b2fc),
	.w5(32'h3b71cdb0),
	.w6(32'h397c707b),
	.w7(32'hb9b31fc5),
	.w8(32'h3b91f6e8),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd7c24a),
	.w1(32'h3b569f95),
	.w2(32'h3b0d88a2),
	.w3(32'h38350ab9),
	.w4(32'h3901e793),
	.w5(32'hb9d679b9),
	.w6(32'h3b5dfa0b),
	.w7(32'h3af59832),
	.w8(32'h3b0173f5),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9d45da),
	.w1(32'h3a9f1ec9),
	.w2(32'h3a43bb44),
	.w3(32'hbb9fc44c),
	.w4(32'hbb567f7d),
	.w5(32'h3a2e397f),
	.w6(32'hbaff12dc),
	.w7(32'hba13ab21),
	.w8(32'hbb734da0),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0071f5),
	.w1(32'h382cc1f6),
	.w2(32'h3ae94678),
	.w3(32'h3ae8cbc1),
	.w4(32'h3b8a909e),
	.w5(32'hbab1d984),
	.w6(32'hbaf73d2b),
	.w7(32'h3a971478),
	.w8(32'hba9c0582),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8ad684),
	.w1(32'hbaeb90a0),
	.w2(32'hba3d074c),
	.w3(32'hbab8af19),
	.w4(32'hb95565f9),
	.w5(32'hbb2b5aaa),
	.w6(32'hbb116a5b),
	.w7(32'hba249da2),
	.w8(32'hbb27ec6d),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9b9e79),
	.w1(32'hbb941fc1),
	.w2(32'hbacc0e7c),
	.w3(32'hbaeb8e3b),
	.w4(32'hba3458e8),
	.w5(32'hb9a4ad73),
	.w6(32'hbb062be2),
	.w7(32'hba48c4dd),
	.w8(32'h3abcb6e6),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4f697e),
	.w1(32'h3b200b54),
	.w2(32'h3a29130a),
	.w3(32'hbb37d4b6),
	.w4(32'h3a3af646),
	.w5(32'h3a73eaef),
	.w6(32'h3aefd7fe),
	.w7(32'h3b1b8f1b),
	.w8(32'h39ae64b2),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7c6b5c),
	.w1(32'h3ac30dfc),
	.w2(32'h3a271f05),
	.w3(32'h3a3ac801),
	.w4(32'h3a994b2f),
	.w5(32'h3b2ac5e0),
	.w6(32'h3b8408f7),
	.w7(32'h3b0e8034),
	.w8(32'h3b86f0eb),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba3804e),
	.w1(32'hb97922a6),
	.w2(32'h3b8146ab),
	.w3(32'hb9a39f67),
	.w4(32'h3b8beb8a),
	.w5(32'hbb060f17),
	.w6(32'h394d3a15),
	.w7(32'h3bb3c315),
	.w8(32'hbb3adc03),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3905c3),
	.w1(32'hba171784),
	.w2(32'hbaee9ead),
	.w3(32'hba4e087d),
	.w4(32'hbb344e68),
	.w5(32'hbb989760),
	.w6(32'hbb2dcc6c),
	.w7(32'hbac7d1d9),
	.w8(32'hbbc2f23b),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbbea8f1),
	.w1(32'hbb6fb340),
	.w2(32'hbb36fa26),
	.w3(32'hbae872df),
	.w4(32'hbae6e53e),
	.w5(32'h3b19febe),
	.w6(32'hbb194430),
	.w7(32'hbb779c4a),
	.w8(32'h3b248076),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3abe88a0),
	.w1(32'h3a8d601b),
	.w2(32'h379778ec),
	.w3(32'hbaf77ca1),
	.w4(32'hbaad52d9),
	.w5(32'hbb984a34),
	.w6(32'h3b28b5f4),
	.w7(32'h38d8cb4c),
	.w8(32'hbbbc91f8),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6ef26a),
	.w1(32'hbab19eab),
	.w2(32'hbb60727f),
	.w3(32'hbaade5e7),
	.w4(32'hbaeb20bd),
	.w5(32'h3b5208bb),
	.w6(32'hbb17f932),
	.w7(32'hbb9da88e),
	.w8(32'h3b2b5591),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a377d36),
	.w1(32'h3a03a5ff),
	.w2(32'h3a0daf54),
	.w3(32'h3b195a38),
	.w4(32'hb75316ed),
	.w5(32'hba8f2e3d),
	.w6(32'h3a5fec38),
	.w7(32'h3a10c844),
	.w8(32'hbacf15ed),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab49366),
	.w1(32'hbb422aec),
	.w2(32'hbb1b7562),
	.w3(32'hbb0bfdb0),
	.w4(32'hbb15da2a),
	.w5(32'hbb099656),
	.w6(32'hbb645bc7),
	.w7(32'hbafe5177),
	.w8(32'hbaf2380b),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8835b65),
	.w1(32'hba62506c),
	.w2(32'hbb098188),
	.w3(32'hbb0879e2),
	.w4(32'hbb26521a),
	.w5(32'h3b924455),
	.w6(32'hbb679ed6),
	.w7(32'hbb50be34),
	.w8(32'h3b0c54b9),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a7ffb11),
	.w1(32'h3a71a4b6),
	.w2(32'hb87f7f7f),
	.w3(32'h3ac048c1),
	.w4(32'h3952fb9a),
	.w5(32'hbafcfde4),
	.w6(32'h3ac2b146),
	.w7(32'h3a7378cd),
	.w8(32'hbad5c1f0),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0e2e54),
	.w1(32'h3c080506),
	.w2(32'h3b0d5389),
	.w3(32'h3be172cd),
	.w4(32'h3b548356),
	.w5(32'h3ae3673b),
	.w6(32'h3c1dddc4),
	.w7(32'hb78d0d93),
	.w8(32'h3b266809),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8ddd327),
	.w1(32'hbb48d927),
	.w2(32'h3b9bed7d),
	.w3(32'hba87cac2),
	.w4(32'hbb818d12),
	.w5(32'h3aaff045),
	.w6(32'h3b0a4f4f),
	.w7(32'h395ffafd),
	.w8(32'h3b45ed95),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1acd67),
	.w1(32'h3bcf7650),
	.w2(32'h3acde7bf),
	.w3(32'h3b7ff0fb),
	.w4(32'h3b608461),
	.w5(32'h3ac183f1),
	.w6(32'h3b8d02d6),
	.w7(32'h3abcdab1),
	.w8(32'h3b520766),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fede20),
	.w1(32'hb8fb732f),
	.w2(32'h3b53f298),
	.w3(32'h3b066807),
	.w4(32'h3a4c55d4),
	.w5(32'hbb945366),
	.w6(32'h3b1fd9c4),
	.w7(32'hba6feb34),
	.w8(32'hbba282b4),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e3f4e),
	.w1(32'hbb7cba9c),
	.w2(32'hbb1f0f6e),
	.w3(32'hb9c3509c),
	.w4(32'hbaf5ab02),
	.w5(32'hbb480380),
	.w6(32'hba752b5a),
	.w7(32'hba1db2e3),
	.w8(32'hbbb59a92),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb98efbb),
	.w1(32'hbb8c755f),
	.w2(32'h3aa5d3c3),
	.w3(32'hb42a1164),
	.w4(32'h3b116c61),
	.w5(32'hb6f25de4),
	.w6(32'hbb79593a),
	.w7(32'hba32fc91),
	.w8(32'hbaa7a452),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeaea9c),
	.w1(32'h3ad63c19),
	.w2(32'h39476a45),
	.w3(32'h3b1efdf0),
	.w4(32'h3af3515f),
	.w5(32'h3b2214c6),
	.w6(32'h3a468443),
	.w7(32'h3ac00c7b),
	.w8(32'h3b847956),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule