module layer_8_featuremap_244(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb0609e7),
	.w1(32'hba1f7ed5),
	.w2(32'h3c2a0f40),
	.w3(32'h3beb1769),
	.w4(32'hba9f3fd0),
	.w5(32'h3d1b8dd4),
	.w6(32'hbbd34e6e),
	.w7(32'hbbb5cefc),
	.w8(32'hbc041246),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb33f1d),
	.w1(32'hbb0c3940),
	.w2(32'hbac25520),
	.w3(32'h3ce45cac),
	.w4(32'hbb3572ae),
	.w5(32'hbb31ece4),
	.w6(32'h3ab4c190),
	.w7(32'h3b088d05),
	.w8(32'h3a7d9481),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7b5466),
	.w1(32'h3b177324),
	.w2(32'h3bc33c5d),
	.w3(32'hba37baa5),
	.w4(32'h3acca5ad),
	.w5(32'hbbdc54a3),
	.w6(32'hba795d3d),
	.w7(32'h3bdd7bc8),
	.w8(32'hbabeb249),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b143447),
	.w1(32'hbb9e6650),
	.w2(32'hbc106203),
	.w3(32'hbbb4dc9d),
	.w4(32'hbbe4d066),
	.w5(32'hbc791a4d),
	.w6(32'h3ad00be3),
	.w7(32'hba87613e),
	.w8(32'hbb793e33),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3f22b6),
	.w1(32'hb7ea950c),
	.w2(32'h39e394ae),
	.w3(32'hbb86431c),
	.w4(32'hbaa79b87),
	.w5(32'h3b0238ac),
	.w6(32'h3b40dde8),
	.w7(32'h39a3bbcd),
	.w8(32'hb9811c48),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b1f372),
	.w1(32'h3b2b6eaa),
	.w2(32'hbc0d3c9f),
	.w3(32'h3b6fafc0),
	.w4(32'hba5b86b3),
	.w5(32'hbc5f013f),
	.w6(32'hbb9450f5),
	.w7(32'hbb47deb5),
	.w8(32'hbacfabc3),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfd5db1),
	.w1(32'hba23e4e8),
	.w2(32'h3a598fb7),
	.w3(32'hbc6f27ec),
	.w4(32'h3b0fdb86),
	.w5(32'h3b7f5600),
	.w6(32'hbb3a882e),
	.w7(32'hbb04f55d),
	.w8(32'hba8048b3),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba22a946),
	.w1(32'h3c488c8f),
	.w2(32'h3baf7520),
	.w3(32'h3b107f21),
	.w4(32'h3b95265b),
	.w5(32'h3b9ad231),
	.w6(32'h3af3c8a2),
	.w7(32'hbbf4011c),
	.w8(32'h3b0e6efe),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bced334),
	.w1(32'hbad0ffa6),
	.w2(32'hbb62a74b),
	.w3(32'hbba64504),
	.w4(32'hbb620127),
	.w5(32'hbba04aa3),
	.w6(32'h3b4a1f8b),
	.w7(32'h3a844151),
	.w8(32'hba20f7e4),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6a6ec5),
	.w1(32'hbba5a7d1),
	.w2(32'hbb6bf030),
	.w3(32'hbb8906a0),
	.w4(32'hba94dc17),
	.w5(32'h3b106365),
	.w6(32'h3be177d4),
	.w7(32'h3b6112ea),
	.w8(32'h3c243bd0),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3dd7f2),
	.w1(32'hb9a53603),
	.w2(32'hbc19331c),
	.w3(32'h3b40afbf),
	.w4(32'hba704315),
	.w5(32'hbc496518),
	.w6(32'hbb02d814),
	.w7(32'hba74846f),
	.w8(32'hbc1a7aae),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba251fa),
	.w1(32'hbb104046),
	.w2(32'hbb0211aa),
	.w3(32'hbc291ed6),
	.w4(32'h3b7351b2),
	.w5(32'h3bad257b),
	.w6(32'hbaa28220),
	.w7(32'hbb2ae856),
	.w8(32'hbb11d750),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaba983b),
	.w1(32'hbab7bc2f),
	.w2(32'hbb3fe2ca),
	.w3(32'h3b80e3f9),
	.w4(32'h3ada64b1),
	.w5(32'hbaddf179),
	.w6(32'h3b941637),
	.w7(32'h3b30a075),
	.w8(32'h3b97be8d),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc09d186),
	.w1(32'hbbad8741),
	.w2(32'hbb062cc2),
	.w3(32'h3b42bb1c),
	.w4(32'hb98781b3),
	.w5(32'hbc1308fd),
	.w6(32'h3adeb689),
	.w7(32'hbae0762f),
	.w8(32'h3bc808a1),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b117439),
	.w1(32'h3b828860),
	.w2(32'h3965892a),
	.w3(32'hbc42fa9c),
	.w4(32'h3b2058c4),
	.w5(32'hbb5c6f9f),
	.w6(32'h3b285c3d),
	.w7(32'h3ada853b),
	.w8(32'h3b03e673),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a00e204),
	.w1(32'hbb9a78b0),
	.w2(32'hbc1dcfb6),
	.w3(32'hbb850f94),
	.w4(32'hbbddbd93),
	.w5(32'h3c8b3420),
	.w6(32'hbb8e121c),
	.w7(32'hbc1c580f),
	.w8(32'hbc1c91e6),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2062e7),
	.w1(32'hbb5f33f9),
	.w2(32'h3be44a09),
	.w3(32'h3cfe342d),
	.w4(32'h3b3c5843),
	.w5(32'h3d44acc3),
	.w6(32'h3c0ae6bf),
	.w7(32'h3b217154),
	.w8(32'hbb82aa5e),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc511cf),
	.w1(32'hbaf7f2d1),
	.w2(32'hbb3b60be),
	.w3(32'h3d4ffe8c),
	.w4(32'h3b12aa83),
	.w5(32'hb9ec9eae),
	.w6(32'h3a5fd51c),
	.w7(32'h3b98fe29),
	.w8(32'h3a0f30f7),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aea2250),
	.w1(32'h3ba017fd),
	.w2(32'h3ab178d8),
	.w3(32'hbb9b55c7),
	.w4(32'hbade3201),
	.w5(32'h3ba918e7),
	.w6(32'h3c126828),
	.w7(32'h3c1aeef2),
	.w8(32'h3c087024),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa7f21b),
	.w1(32'h39386dc4),
	.w2(32'hbad8a0fd),
	.w3(32'hbbe7da31),
	.w4(32'hb7623785),
	.w5(32'hbba55e44),
	.w6(32'hb9d84ee9),
	.w7(32'hba140a47),
	.w8(32'hb9c5d3be),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac41804),
	.w1(32'hbb2d6499),
	.w2(32'h3c1925a2),
	.w3(32'hbb8c28e4),
	.w4(32'h3beb47dd),
	.w5(32'h3d0d7ea1),
	.w6(32'h3a4d7963),
	.w7(32'hbc18d7fc),
	.w8(32'hbbecd21b),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb00c1e6),
	.w1(32'h3c7e94d4),
	.w2(32'h3ab40c33),
	.w3(32'h3cacf08c),
	.w4(32'hbb863638),
	.w5(32'hbc587ab4),
	.w6(32'h3966d5c4),
	.w7(32'hbb09c367),
	.w8(32'h3ae691de),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9a5712),
	.w1(32'h3b952a61),
	.w2(32'hbb79a8f2),
	.w3(32'hbb430373),
	.w4(32'hbc1593c2),
	.w5(32'hbc5b37ba),
	.w6(32'h3bdd6935),
	.w7(32'h3bc39251),
	.w8(32'h3bd74498),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba5a5d8),
	.w1(32'h3bd4e971),
	.w2(32'h3b368ed1),
	.w3(32'hbb280700),
	.w4(32'hbb35a8ad),
	.w5(32'hb897a760),
	.w6(32'h391b223a),
	.w7(32'hbb4a40e7),
	.w8(32'hbb69fe91),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbac3d73),
	.w1(32'h39132c31),
	.w2(32'hba59c12d),
	.w3(32'hbbb4ad64),
	.w4(32'h3a2b6105),
	.w5(32'hbb02ce06),
	.w6(32'h3a834195),
	.w7(32'hbaf42b9c),
	.w8(32'hb9b38e56),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1647c3),
	.w1(32'hba2d4856),
	.w2(32'h3cb3578f),
	.w3(32'h3aa0dcd6),
	.w4(32'hbba88287),
	.w5(32'h3bd30dff),
	.w6(32'hbc279949),
	.w7(32'hbaae504c),
	.w8(32'hbb8614e7),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8d6845),
	.w1(32'h3a61abf2),
	.w2(32'hbb25d76c),
	.w3(32'h3b12b6fd),
	.w4(32'hbc0e877c),
	.w5(32'hbc016918),
	.w6(32'hbae93444),
	.w7(32'hba591097),
	.w8(32'hbb049039),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8a0f58),
	.w1(32'hbb77cd37),
	.w2(32'hbbe2badf),
	.w3(32'hbba8a21d),
	.w4(32'hbc05b495),
	.w5(32'hbc526760),
	.w6(32'h3926ca25),
	.w7(32'hb983adfc),
	.w8(32'hbc0edd37),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba85ba0d),
	.w1(32'hbae48163),
	.w2(32'h3b8be857),
	.w3(32'hbc0bfdd9),
	.w4(32'hbaf25248),
	.w5(32'h3b398f26),
	.w6(32'hbbaa38dd),
	.w7(32'hb86cb5e0),
	.w8(32'hbac5343c),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9c4749),
	.w1(32'hba41d501),
	.w2(32'hb9a7bd12),
	.w3(32'hbc0460ad),
	.w4(32'h3bb83ed3),
	.w5(32'h3b923d8a),
	.w6(32'hba46ad1e),
	.w7(32'hbae3d10d),
	.w8(32'hbbc808ed),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb2b1f0),
	.w1(32'h3b0cd54e),
	.w2(32'h3c008bac),
	.w3(32'h39093b64),
	.w4(32'h39a23110),
	.w5(32'h3ba4cb8c),
	.w6(32'hbb722e5f),
	.w7(32'h3a29f33c),
	.w8(32'hbb2f0515),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0436be),
	.w1(32'hbb34cdda),
	.w2(32'h3b9bc54d),
	.w3(32'h3b9e75a9),
	.w4(32'h3a46200e),
	.w5(32'h3c68c17f),
	.w6(32'hba8b80c5),
	.w7(32'hba40ffa4),
	.w8(32'hbaa69416),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9a6182),
	.w1(32'hba7e192c),
	.w2(32'hba9ccde4),
	.w3(32'h3cb4d80f),
	.w4(32'h3ba672ed),
	.w5(32'hbc203a90),
	.w6(32'h3bce6436),
	.w7(32'h3b9c3206),
	.w8(32'hb7e4a604),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1136fa),
	.w1(32'h3a7cc1c2),
	.w2(32'h3bc64c90),
	.w3(32'hbba2fc45),
	.w4(32'hbaf065c5),
	.w5(32'h3c05a476),
	.w6(32'h3af243c7),
	.w7(32'hba5be26c),
	.w8(32'hbbcca44a),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b25a2f8),
	.w1(32'h3a93c21b),
	.w2(32'hbb48ee87),
	.w3(32'h3b2217a4),
	.w4(32'h3b125d7e),
	.w5(32'h3b1b651f),
	.w6(32'h3b3811f5),
	.w7(32'h3a971036),
	.w8(32'hb938324a),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3985a672),
	.w1(32'h3b1a2b0d),
	.w2(32'h3ba4da45),
	.w3(32'h3b4bdb62),
	.w4(32'h3a7197d5),
	.w5(32'h3b955291),
	.w6(32'hba48c866),
	.w7(32'h3b27a251),
	.w8(32'hbb6edaa7),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b90c3cd),
	.w1(32'h3956812e),
	.w2(32'h3b17a1e9),
	.w3(32'hbaea0f5e),
	.w4(32'hb99b9ccb),
	.w5(32'h39821249),
	.w6(32'h3a54db79),
	.w7(32'h3aab4348),
	.w8(32'hb9b84f52),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37cbfe80),
	.w1(32'h3b4a1a9a),
	.w2(32'hbb51e8fe),
	.w3(32'hbabb6400),
	.w4(32'h3a401dc2),
	.w5(32'hbbe0554a),
	.w6(32'h3bbdcdf3),
	.w7(32'h3aea1349),
	.w8(32'h3a98f2dc),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb25aa36),
	.w1(32'h3b016970),
	.w2(32'hbb34cec1),
	.w3(32'hbbb9c13d),
	.w4(32'hbab85a1a),
	.w5(32'hbb2698c3),
	.w6(32'hbafc5df1),
	.w7(32'hbb7e2061),
	.w8(32'h3aaff799),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc086c21),
	.w1(32'h3bab1c06),
	.w2(32'h3b446c7d),
	.w3(32'hbbbc4f07),
	.w4(32'hbb69942e),
	.w5(32'h3b593d02),
	.w6(32'hba7088e6),
	.w7(32'hbb99c2d5),
	.w8(32'hbbb6b5d9),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2b6586),
	.w1(32'hb9ba53bb),
	.w2(32'h39766f31),
	.w3(32'h3af8eaad),
	.w4(32'hb85cf5b4),
	.w5(32'hba8439e6),
	.w6(32'h391e7c31),
	.w7(32'h3a3fc0ae),
	.w8(32'h38d9c05a),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h381da97f),
	.w1(32'hba83cab9),
	.w2(32'hba83b3ea),
	.w3(32'hba9ee054),
	.w4(32'h3a8eb7a8),
	.w5(32'hbaf3e5de),
	.w6(32'hbae76af6),
	.w7(32'hbb88b04d),
	.w8(32'hbb8bbe0f),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc89e13),
	.w1(32'hbb253ee2),
	.w2(32'h3b0e72c3),
	.w3(32'h3bf5e35a),
	.w4(32'h3a98054e),
	.w5(32'hb98e4043),
	.w6(32'hba90b2ff),
	.w7(32'h3b05971a),
	.w8(32'hba15402e),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39de7dd7),
	.w1(32'hbba7db98),
	.w2(32'hbbbf66b6),
	.w3(32'h3b815ce9),
	.w4(32'h3c27bb51),
	.w5(32'h3a1393b9),
	.w6(32'h3b8330cd),
	.w7(32'h3b63ba87),
	.w8(32'hbac34ac2),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9695db),
	.w1(32'hbab2af43),
	.w2(32'h3b20d577),
	.w3(32'h3b19e219),
	.w4(32'hbcaa2b90),
	.w5(32'hbce2a8fc),
	.w6(32'h3bc16854),
	.w7(32'h3ba4a59a),
	.w8(32'hb9ecbe7a),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2171d2),
	.w1(32'hba9bf541),
	.w2(32'h3a78b838),
	.w3(32'hbca72a77),
	.w4(32'hbaa56881),
	.w5(32'hba805d68),
	.w6(32'hbaddec6e),
	.w7(32'hba19ff9f),
	.w8(32'hbaf34612),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba62dffd),
	.w1(32'hba9d957e),
	.w2(32'h3bb3ae9a),
	.w3(32'hbb1ab505),
	.w4(32'h396da812),
	.w5(32'h3c0c6c40),
	.w6(32'hbb7de7d1),
	.w7(32'hbb0cbc7c),
	.w8(32'h3b0991a4),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf7fceb),
	.w1(32'h3b91fcdf),
	.w2(32'hb9942180),
	.w3(32'h3c6fbb4f),
	.w4(32'h3b4966c0),
	.w5(32'hbba6a086),
	.w6(32'h3b848c48),
	.w7(32'hbae5c3c7),
	.w8(32'hbb836d98),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb61edb8),
	.w1(32'h3c086609),
	.w2(32'h3b2591a6),
	.w3(32'hbb06e8ac),
	.w4(32'hbb4a604d),
	.w5(32'hbbeb5517),
	.w6(32'h3c2390ad),
	.w7(32'hbaea2133),
	.w8(32'h3add4ae6),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2c883c),
	.w1(32'hbb1f3c64),
	.w2(32'hbaa04a02),
	.w3(32'h3b18a7cd),
	.w4(32'hbaa4463c),
	.w5(32'hbc3af0da),
	.w6(32'h3bd820a0),
	.w7(32'h3a5fc5cf),
	.w8(32'h3ae7fd3f),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1da10a),
	.w1(32'hba000e5e),
	.w2(32'h3a396cdd),
	.w3(32'hbae139ff),
	.w4(32'h37a5848d),
	.w5(32'h3a95fe6d),
	.w6(32'hba2697c4),
	.w7(32'h3af6aec0),
	.w8(32'hba957567),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba636407),
	.w1(32'h3a8e9e0c),
	.w2(32'h3a188783),
	.w3(32'hba1e4eab),
	.w4(32'hba3ffde5),
	.w5(32'hba3da640),
	.w6(32'hbb15e975),
	.w7(32'h3aaff4b9),
	.w8(32'hba86e7cf),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaedcbe7),
	.w1(32'hba47e232),
	.w2(32'hbb357466),
	.w3(32'hba946dcd),
	.w4(32'hba727fb3),
	.w5(32'hbad82880),
	.w6(32'h3b35cddd),
	.w7(32'h3a4702c4),
	.w8(32'hba4f72c8),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb88b92e),
	.w1(32'hbc0844b3),
	.w2(32'h3b25d214),
	.w3(32'hbaa1468c),
	.w4(32'h3cc7ad09),
	.w5(32'h3d23a4f3),
	.w6(32'hbc44cee0),
	.w7(32'hbc71f8dd),
	.w8(32'hbbc85d7b),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h37edc000),
	.w1(32'hbb24f1ae),
	.w2(32'hbc0a5183),
	.w3(32'h3c887d19),
	.w4(32'hbb3f2121),
	.w5(32'hbc652a8f),
	.w6(32'h3c0df69d),
	.w7(32'h3b10a487),
	.w8(32'hba35b159),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc477340),
	.w1(32'hbbad7310),
	.w2(32'hbc0cd6ba),
	.w3(32'hbc1eadfe),
	.w4(32'h3be91be4),
	.w5(32'hba625d0f),
	.w6(32'h398a0bf1),
	.w7(32'h3b518b27),
	.w8(32'hbb2c9bb7),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b36b384),
	.w1(32'h39bcc69f),
	.w2(32'hbc128b92),
	.w3(32'hbbd39ede),
	.w4(32'hbb1a9309),
	.w5(32'hbc7f7deb),
	.w6(32'h3bda81bd),
	.w7(32'h3b5fb4b2),
	.w8(32'hb9e64b37),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb849c7a),
	.w1(32'h3a05f2fe),
	.w2(32'h3b4d65f4),
	.w3(32'hbaa4df71),
	.w4(32'h3b78337e),
	.w5(32'h3b9e323a),
	.w6(32'hba66c995),
	.w7(32'h3b679b3d),
	.w8(32'h3ab31f0c),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b01dafc),
	.w1(32'hbab38c4e),
	.w2(32'h394ddda1),
	.w3(32'hb8b69690),
	.w4(32'hbaccd41f),
	.w5(32'hba9a73d1),
	.w6(32'h3a8db7c5),
	.w7(32'h39cb2d07),
	.w8(32'h3b3d1930),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b274e7a),
	.w1(32'h3c2938f6),
	.w2(32'h3c16f82e),
	.w3(32'h3ac8404f),
	.w4(32'hb8d1b408),
	.w5(32'hbbf0609c),
	.w6(32'h3b4f5a91),
	.w7(32'hbb6f8d23),
	.w8(32'h37fe64d2),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9d494e),
	.w1(32'hbbcefd67),
	.w2(32'hbc35c310),
	.w3(32'h3aad8ca2),
	.w4(32'hbb82f54b),
	.w5(32'hbc4732ec),
	.w6(32'hba693802),
	.w7(32'hbb0907a8),
	.w8(32'h3a0128b7),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba37c4f),
	.w1(32'hbb91f2f5),
	.w2(32'hba1b0ab0),
	.w3(32'h39eba22d),
	.w4(32'hbb8acd4f),
	.w5(32'hb8df3077),
	.w6(32'hbb1b5eff),
	.w7(32'hbb7c85ff),
	.w8(32'hba2c38c6),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb044725),
	.w1(32'hbb7a736f),
	.w2(32'hbb11ced5),
	.w3(32'h3aec9c17),
	.w4(32'hbaee6b80),
	.w5(32'h3bddd215),
	.w6(32'hba8fd080),
	.w7(32'hbaa82d60),
	.w8(32'hb7c89b6c),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd991a8),
	.w1(32'hbb950ac2),
	.w2(32'hbc15e711),
	.w3(32'h3b999ba7),
	.w4(32'hbb1c8537),
	.w5(32'hbb9f14cf),
	.w6(32'hbb65b6cc),
	.w7(32'hbb495154),
	.w8(32'hbb2de0d5),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb9adb3),
	.w1(32'h39274c5b),
	.w2(32'hba54312d),
	.w3(32'hba0ea48f),
	.w4(32'hb9541bb3),
	.w5(32'hba8a6553),
	.w6(32'h39d3ac53),
	.w7(32'h3a892cc2),
	.w8(32'h3ab5ec7c),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba0a15e3),
	.w1(32'h3acab0b6),
	.w2(32'h3abd0a0d),
	.w3(32'hbb060783),
	.w4(32'h3aea27e9),
	.w5(32'h3bb40877),
	.w6(32'hbafd368f),
	.w7(32'hbbac7204),
	.w8(32'h3adb8b1d),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba89504),
	.w1(32'hbbf833fe),
	.w2(32'hbbec8cdb),
	.w3(32'h3b957650),
	.w4(32'hbaa55725),
	.w5(32'h3cc03909),
	.w6(32'h3a4c1687),
	.w7(32'hbbc3e4c9),
	.w8(32'hbbba43be),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc20f8bb),
	.w1(32'hbc4281d6),
	.w2(32'hba401d34),
	.w3(32'h3ce37107),
	.w4(32'hbbdfa775),
	.w5(32'hb871af1c),
	.w6(32'hbc1b5c43),
	.w7(32'hbc6490df),
	.w8(32'hbc50306b),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbaccf8e),
	.w1(32'hbbf033c8),
	.w2(32'hbb3b8f94),
	.w3(32'hbba0ee07),
	.w4(32'hbb2ff648),
	.w5(32'hbaa712f7),
	.w6(32'hbb668dc1),
	.w7(32'hbae8d5f1),
	.w8(32'h39d2cb84),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baa0090),
	.w1(32'h3be4cc37),
	.w2(32'h3b2e82d1),
	.w3(32'hba4a7307),
	.w4(32'hbb321ae3),
	.w5(32'hbbd3e2ed),
	.w6(32'h3adb0b3b),
	.w7(32'h3bc9817b),
	.w8(32'h3bbfbb5a),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb695c77),
	.w1(32'hbb0ec0de),
	.w2(32'hbbb03958),
	.w3(32'h3b619d87),
	.w4(32'h3a99b90a),
	.w5(32'hba0ab2f4),
	.w6(32'hbba08718),
	.w7(32'hbbd85fe6),
	.w8(32'hbb194996),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9693f2a),
	.w1(32'hba6fd938),
	.w2(32'h3c04b609),
	.w3(32'h3b7eb6fc),
	.w4(32'hbb9265a6),
	.w5(32'hba1c5549),
	.w6(32'hbb99be0b),
	.w7(32'h3bdd2062),
	.w8(32'h3b13f97d),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8acb86),
	.w1(32'h3a27eff7),
	.w2(32'h395b808b),
	.w3(32'hbb68322e),
	.w4(32'hbac7d68a),
	.w5(32'hbb8f54e1),
	.w6(32'h3b33ebe1),
	.w7(32'h3ba195a5),
	.w8(32'h3b31339e),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bfd9a4f),
	.w1(32'h3a692699),
	.w2(32'hbac33360),
	.w3(32'hbb52ce05),
	.w4(32'h3a37b5bf),
	.w5(32'hbb0e4e2a),
	.w6(32'h3ad964e3),
	.w7(32'h3a8a301e),
	.w8(32'h3a761707),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbeb9fb),
	.w1(32'hb900f5d9),
	.w2(32'hb98c3c23),
	.w3(32'h3af60079),
	.w4(32'hbb7d297b),
	.w5(32'hbabecf6f),
	.w6(32'h3ae0dea2),
	.w7(32'h3b11b27e),
	.w8(32'hb9e481ba),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b21e79a),
	.w1(32'h3bc5a540),
	.w2(32'h39c42d27),
	.w3(32'h3a3f458c),
	.w4(32'h3ba0d166),
	.w5(32'hbad31e46),
	.w6(32'h3c05fcf2),
	.w7(32'h3c16cb5d),
	.w8(32'h3be7cc90),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a43daf5),
	.w1(32'h3b41a6f6),
	.w2(32'h3b0d7bf3),
	.w3(32'h3c514b9f),
	.w4(32'h3bcbe5cd),
	.w5(32'h3bd02a5d),
	.w6(32'hba866c6a),
	.w7(32'h3acad4ba),
	.w8(32'h3b56a585),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa099f3),
	.w1(32'hbb00e2dd),
	.w2(32'h3a811397),
	.w3(32'h3bc85d40),
	.w4(32'hbac920e3),
	.w5(32'hbacdac5e),
	.w6(32'hba97f463),
	.w7(32'h3b80289a),
	.w8(32'hb7829e6f),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aaac9bb),
	.w1(32'hbb131c92),
	.w2(32'hbb3b1eb3),
	.w3(32'h39335992),
	.w4(32'h3bf0a62e),
	.w5(32'h3985725d),
	.w6(32'hbba3a6f4),
	.w7(32'h3ac26703),
	.w8(32'h3b91cd0f),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9fa66ed),
	.w1(32'hbc193e6f),
	.w2(32'hbb0c0417),
	.w3(32'hba9c69df),
	.w4(32'hbab518b0),
	.w5(32'h3ba30057),
	.w6(32'h39c06da6),
	.w7(32'hbb0b2791),
	.w8(32'h3aae6573),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c290ba1),
	.w1(32'hb96146e7),
	.w2(32'h3b8d437f),
	.w3(32'h3b956016),
	.w4(32'h3b054738),
	.w5(32'hb90c43c1),
	.w6(32'hba293ec4),
	.w7(32'h3b2b92af),
	.w8(32'h3b32793d),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf06454),
	.w1(32'hbb4431b6),
	.w2(32'h3bb78608),
	.w3(32'hbb62bc07),
	.w4(32'hba1f72d7),
	.w5(32'hba05f7ab),
	.w6(32'hbba96377),
	.w7(32'hbb882466),
	.w8(32'hbb36afb7),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baa181d),
	.w1(32'h3b92700f),
	.w2(32'hbb58fec6),
	.w3(32'hbbcc89ef),
	.w4(32'h3a6e8071),
	.w5(32'hbbe049d2),
	.w6(32'h3ba00b98),
	.w7(32'h3c00baca),
	.w8(32'h3b3d39b0),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb84f7db),
	.w1(32'hbc1be22a),
	.w2(32'hbba52125),
	.w3(32'hba9823cf),
	.w4(32'hb8f13af9),
	.w5(32'h3addada5),
	.w6(32'hbb8436e7),
	.w7(32'hbbbfa353),
	.w8(32'hbc0291ca),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0ce095),
	.w1(32'h3b0629e1),
	.w2(32'h3aa7eead),
	.w3(32'hbbf22505),
	.w4(32'hbb9c24b8),
	.w5(32'hbc269d23),
	.w6(32'h3bb0d2d4),
	.w7(32'h3be6cac5),
	.w8(32'h3b45c481),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ab42332),
	.w1(32'hbb1c62d7),
	.w2(32'hbc2e0f46),
	.w3(32'hbc0175d7),
	.w4(32'hbbcbc196),
	.w5(32'hbb6c0627),
	.w6(32'hbc06ea55),
	.w7(32'hba4d9530),
	.w8(32'hbb8b8bff),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe36680),
	.w1(32'hbb80457f),
	.w2(32'hb9521f69),
	.w3(32'hbb2b0bbb),
	.w4(32'hbbd742b7),
	.w5(32'hbbb20baf),
	.w6(32'hbb2cec6f),
	.w7(32'hbacf3dce),
	.w8(32'hbac0d41e),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa4e92e),
	.w1(32'hbba21066),
	.w2(32'hbc028657),
	.w3(32'hbba8a238),
	.w4(32'h3b4079d7),
	.w5(32'h3a8273d1),
	.w6(32'h3b54c2c1),
	.w7(32'h39c7d050),
	.w8(32'h3bcd760c),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf43911),
	.w1(32'hb9c28d14),
	.w2(32'h3b2a4d87),
	.w3(32'h3abc24c6),
	.w4(32'hba842acf),
	.w5(32'h39fd7287),
	.w6(32'hbb389f40),
	.w7(32'hbb05ef4b),
	.w8(32'hbb8c1d3c),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac928ae),
	.w1(32'h3aaf08e6),
	.w2(32'h3b9dbb38),
	.w3(32'h3a06180f),
	.w4(32'hb9d665f3),
	.w5(32'hbc85f25b),
	.w6(32'h3be24dcf),
	.w7(32'h3a564bc3),
	.w8(32'hbb48a07e),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba3d20e),
	.w1(32'hbb643eb6),
	.w2(32'h3bc6e3a5),
	.w3(32'hbc37f5df),
	.w4(32'hbb957bb4),
	.w5(32'h39dbdf0f),
	.w6(32'h3c0157b7),
	.w7(32'h3bcd4b01),
	.w8(32'h3a37fb64),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb8a634),
	.w1(32'hbada7b91),
	.w2(32'h3a7c828d),
	.w3(32'hbbc01780),
	.w4(32'hbb61629e),
	.w5(32'h3c61a227),
	.w6(32'hbb4ac8fe),
	.w7(32'hbaaec97f),
	.w8(32'hbb5bcf04),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba212343),
	.w1(32'hbb2da8b0),
	.w2(32'hbba0f4f7),
	.w3(32'h3be5dafe),
	.w4(32'hbb12e54c),
	.w5(32'hbb576106),
	.w6(32'hbae5bd65),
	.w7(32'hbb34d059),
	.w8(32'hbacd5771),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2ed87c),
	.w1(32'hbb18365f),
	.w2(32'hba9873fd),
	.w3(32'h3a70b551),
	.w4(32'hbad9c2eb),
	.w5(32'hba7abe1f),
	.w6(32'hb9aad534),
	.w7(32'hba1f8fab),
	.w8(32'h3870f505),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a6081cd),
	.w1(32'hbab238b1),
	.w2(32'hbba8c523),
	.w3(32'h3b0f7acc),
	.w4(32'hbc2fd6ce),
	.w5(32'hbc164aa9),
	.w6(32'h394a19d4),
	.w7(32'h3bc41e15),
	.w8(32'hbb52038b),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc49c0f),
	.w1(32'hbae56bad),
	.w2(32'hb9d5e9f9),
	.w3(32'hbba342ba),
	.w4(32'hb9a0a4b2),
	.w5(32'h3af7e0ce),
	.w6(32'hbaef61f0),
	.w7(32'hba917665),
	.w8(32'hbba36372),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9e6211),
	.w1(32'h3b9642b1),
	.w2(32'h3bdc6350),
	.w3(32'hbb0bafcb),
	.w4(32'hbbc60ee5),
	.w5(32'hbc07a030),
	.w6(32'h3b5d6556),
	.w7(32'h3b40469d),
	.w8(32'h3b98dcfd),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb17aaa),
	.w1(32'h3a4dcb6c),
	.w2(32'hbba3306b),
	.w3(32'hbc708013),
	.w4(32'h3bd34cb8),
	.w5(32'hbbb1d35e),
	.w6(32'h39500230),
	.w7(32'h3b7af51d),
	.w8(32'h3b83fc08),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1be558),
	.w1(32'h38f059b0),
	.w2(32'hbbc81cb5),
	.w3(32'hbb9e14b9),
	.w4(32'h3c427ead),
	.w5(32'hb927a947),
	.w6(32'hbb753ace),
	.w7(32'hba66a1f6),
	.w8(32'h3a5ad969),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0ff24c),
	.w1(32'h3b7e730c),
	.w2(32'h3b09e0fb),
	.w3(32'h3bde2929),
	.w4(32'h3ae983a4),
	.w5(32'hbbfc9d82),
	.w6(32'h3b5d4ffe),
	.w7(32'h3b0cf596),
	.w8(32'hba051a46),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b5e0f31),
	.w1(32'hba85f4ad),
	.w2(32'h3a9c027b),
	.w3(32'hbabcc632),
	.w4(32'h3c0b5d71),
	.w5(32'h3ccd2c6a),
	.w6(32'hbba7a795),
	.w7(32'hbbdb5c1e),
	.w8(32'hbaba9973),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2171bb),
	.w1(32'hbc4054a3),
	.w2(32'hbc966904),
	.w3(32'hbb1ade82),
	.w4(32'hbc771491),
	.w5(32'hbca7c861),
	.w6(32'h3a018c0a),
	.w7(32'hbb935198),
	.w8(32'hb9d72ccf),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc084583),
	.w1(32'hba3e09ae),
	.w2(32'h3ba66d32),
	.w3(32'hbc78050b),
	.w4(32'hbb99628a),
	.w5(32'h3b6033c8),
	.w6(32'hbad379ce),
	.w7(32'h3b6bb8da),
	.w8(32'h3a9e9754),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6a17e9),
	.w1(32'hbacd49dc),
	.w2(32'hbc4b6a15),
	.w3(32'hbadb8567),
	.w4(32'hbc6584cd),
	.w5(32'hbc6c61cf),
	.w6(32'h3bcde8e5),
	.w7(32'h3ae1d88e),
	.w8(32'hbb9a750e),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc390caf),
	.w1(32'hbb949427),
	.w2(32'hbc475222),
	.w3(32'hbc25d93e),
	.w4(32'h3b08a6ec),
	.w5(32'hbab2699a),
	.w6(32'hbb26d967),
	.w7(32'h3b05075c),
	.w8(32'h3b897b7f),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf93a5b),
	.w1(32'hbada57a3),
	.w2(32'hb8d3c671),
	.w3(32'h3c116dfb),
	.w4(32'hbb0a7c2f),
	.w5(32'h39b6c32a),
	.w6(32'hb9e2792f),
	.w7(32'hb89a0cf7),
	.w8(32'hbacb343a),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb05f32b),
	.w1(32'h37fd1732),
	.w2(32'hbb9f2e67),
	.w3(32'hbb509e91),
	.w4(32'hbbef17a9),
	.w5(32'hba609dac),
	.w6(32'h3b1609de),
	.w7(32'h3b526cad),
	.w8(32'hb913831c),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb981a6d4),
	.w1(32'hba33ce89),
	.w2(32'h3a8449dd),
	.w3(32'h3c1b0a5b),
	.w4(32'h38ef1882),
	.w5(32'hbbbf9b16),
	.w6(32'hbb08cc1e),
	.w7(32'hbac9b9dc),
	.w8(32'hba8deb44),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2ff03a),
	.w1(32'hb6982759),
	.w2(32'h3bad579c),
	.w3(32'h3b3ccf29),
	.w4(32'h3b93cab3),
	.w5(32'h3c9d8246),
	.w6(32'h3b187b54),
	.w7(32'hbaa954a3),
	.w8(32'hbaa1b256),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2ebe12),
	.w1(32'h390491c5),
	.w2(32'h3ab769b4),
	.w3(32'h3c290d76),
	.w4(32'h3a01f932),
	.w5(32'h3b886ebe),
	.w6(32'h3acdaa1c),
	.w7(32'h3a7d9ad0),
	.w8(32'h39c1391b),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391669ca),
	.w1(32'h3a976b19),
	.w2(32'h3b2995e9),
	.w3(32'h3b264701),
	.w4(32'h3a42e3b4),
	.w5(32'h3b426fed),
	.w6(32'hbb485685),
	.w7(32'h3ba1b503),
	.w8(32'hbb608d0f),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3baf6dd1),
	.w1(32'hbb054e6f),
	.w2(32'hb9f2ceb6),
	.w3(32'hb9eff7d7),
	.w4(32'hba39c503),
	.w5(32'hbab41f11),
	.w6(32'hbaab38b8),
	.w7(32'hbabc636c),
	.w8(32'hb9bf1046),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac47795),
	.w1(32'hbbec59c5),
	.w2(32'hbba82524),
	.w3(32'hbaa8bea6),
	.w4(32'hbba585a2),
	.w5(32'hbb8d9377),
	.w6(32'hbbf145f2),
	.w7(32'hbc018278),
	.w8(32'hbaec24f9),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7a9d21),
	.w1(32'hbaead0d7),
	.w2(32'h3a9b5d4d),
	.w3(32'hba625bb0),
	.w4(32'hbba6acd6),
	.w5(32'hbbb70cd0),
	.w6(32'hba9ef275),
	.w7(32'h3af7ac40),
	.w8(32'h3a0f0550),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc05a316),
	.w1(32'h39bace4a),
	.w2(32'h3ae879b1),
	.w3(32'h394eceeb),
	.w4(32'h3a301129),
	.w5(32'h39bf87b6),
	.w6(32'hbad7fcc9),
	.w7(32'h39ca26a8),
	.w8(32'h39e0086a),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0c800d),
	.w1(32'h3ac28139),
	.w2(32'h3aa05e56),
	.w3(32'h3b6b5491),
	.w4(32'h3b1c555c),
	.w5(32'h3aca42c2),
	.w6(32'h3b4011b2),
	.w7(32'h3b75a0a5),
	.w8(32'h3b64f228),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2df2e6),
	.w1(32'hba3fbf79),
	.w2(32'h3b1226ed),
	.w3(32'h3aca297f),
	.w4(32'h3ab78640),
	.w5(32'h3a61d979),
	.w6(32'hba73419c),
	.w7(32'h3b52486b),
	.w8(32'h3acf8bc9),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a169af8),
	.w1(32'h3b141edd),
	.w2(32'h3a0157d3),
	.w3(32'hb9b89b91),
	.w4(32'hbb34adf4),
	.w5(32'hbb6190f4),
	.w6(32'hbb2de085),
	.w7(32'hbb5b3748),
	.w8(32'h3b231faf),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbda2a97),
	.w1(32'hbaa1ed1f),
	.w2(32'hbbf0827a),
	.w3(32'h3a705906),
	.w4(32'h3a2bb7b7),
	.w5(32'hbc686ee7),
	.w6(32'hba19f99b),
	.w7(32'h3a98780b),
	.w8(32'hbacb951b),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc01593e),
	.w1(32'hbb155743),
	.w2(32'hbaba6496),
	.w3(32'hbca82ee2),
	.w4(32'hbb20da1d),
	.w5(32'hbab858ca),
	.w6(32'h3aa83158),
	.w7(32'h3a9bb245),
	.w8(32'hb9b18fe4),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaad6f5e),
	.w1(32'hbbdf1e89),
	.w2(32'h3b8fd250),
	.w3(32'hbb2417cc),
	.w4(32'h3b49df5c),
	.w5(32'h3b7c2376),
	.w6(32'h3b39bef8),
	.w7(32'hbb450439),
	.w8(32'hbb3ee17e),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b1ba2e4),
	.w1(32'h3bc13e4c),
	.w2(32'hbb2d0dcc),
	.w3(32'hbb2c1e37),
	.w4(32'h3b5bb338),
	.w5(32'hbbeba975),
	.w6(32'h3c0c6e28),
	.w7(32'h3bc81c92),
	.w8(32'h3bb79520),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h394e1ac9),
	.w1(32'hbbc8dfaf),
	.w2(32'hbb8d6c11),
	.w3(32'hbc196dd3),
	.w4(32'hbb7094ed),
	.w5(32'hba23a29c),
	.w6(32'hbb30b3e8),
	.w7(32'hbb22ffd6),
	.w8(32'hbb428148),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb38889c),
	.w1(32'h391efcf7),
	.w2(32'hbb0e61ff),
	.w3(32'h391a3f4d),
	.w4(32'hbbb95498),
	.w5(32'hba9ffe12),
	.w6(32'hbb112bbd),
	.w7(32'hbbb3a15b),
	.w8(32'h3954503f),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc135c01),
	.w1(32'hbbad0a3e),
	.w2(32'hbb80dad2),
	.w3(32'h3a901af9),
	.w4(32'h3c3f5a63),
	.w5(32'h3c852d11),
	.w6(32'hbb637b31),
	.w7(32'h3a46373f),
	.w8(32'h3a943efc),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb70f7ed),
	.w1(32'h3c2392a3),
	.w2(32'hb8b38867),
	.w3(32'h3c0f24fb),
	.w4(32'hbbaa4b61),
	.w5(32'hbc04545b),
	.w6(32'h3c07f82a),
	.w7(32'hba5639f2),
	.w8(32'hbafcfe2a),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f9867),
	.w1(32'hbaf692cb),
	.w2(32'hbb8e80ff),
	.w3(32'hbb8f8c5d),
	.w4(32'hbaede790),
	.w5(32'hbb4dd8b6),
	.w6(32'hbb0a2a5c),
	.w7(32'hbb5c66b0),
	.w8(32'hba786dca),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb31c946),
	.w1(32'h3a8d4d63),
	.w2(32'hbb38b414),
	.w3(32'hbaad2961),
	.w4(32'h3b5626e7),
	.w5(32'h3bd1353a),
	.w6(32'hbabed47d),
	.w7(32'hbbc0605d),
	.w8(32'hbc1a7877),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule