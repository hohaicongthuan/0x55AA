module layer_10_featuremap_282(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 8192;
	parameter IMG_SIZE = 13;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc4dfb2),
	.w1(32'hbc11b05a),
	.w2(32'h3cd56ddb),
	.w3(32'hbc4d4f5c),
	.w4(32'h3cbf92d9),
	.w5(32'hbc4cafcc),
	.w6(32'hbd1a1968),
	.w7(32'h3c90f606),
	.w8(32'hbb5f2707),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39a950bd),
	.w1(32'hbb4e6ebc),
	.w2(32'hbc4920ea),
	.w3(32'hbb518b89),
	.w4(32'h3ad5a3f9),
	.w5(32'h3ae36d12),
	.w6(32'hbc3a2c67),
	.w7(32'hbb5266ef),
	.w8(32'h3bad3b29),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1e2a70),
	.w1(32'h3b4064f9),
	.w2(32'hb9bf6d91),
	.w3(32'h3ae68db6),
	.w4(32'hbb3e6cd2),
	.w5(32'hbba7eca2),
	.w6(32'h3c157e56),
	.w7(32'hba7395af),
	.w8(32'h39b27ae1),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba1fefb5),
	.w1(32'h3b65dadf),
	.w2(32'hbbd4a3da),
	.w3(32'h3b43eb95),
	.w4(32'hba2adf54),
	.w5(32'hba8bc0ca),
	.w6(32'h3c6e977a),
	.w7(32'h3b77c4e7),
	.w8(32'hbaee130d),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bc544d3),
	.w1(32'h3c10fb11),
	.w2(32'h3ca708d6),
	.w3(32'h3b72438c),
	.w4(32'h3c6229c3),
	.w5(32'h3b38105f),
	.w6(32'hbb23e2ad),
	.w7(32'h3c90047d),
	.w8(32'hbb8725e9),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h36f0426f),
	.w1(32'hbc0cbf0b),
	.w2(32'hba878405),
	.w3(32'hbba95fa3),
	.w4(32'h3b11219b),
	.w5(32'hb9e94770),
	.w6(32'hbc8d224e),
	.w7(32'hbbc261ac),
	.w8(32'hba6b4928),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a209f52),
	.w1(32'hbc204ec3),
	.w2(32'hbc28b44b),
	.w3(32'hb94696cd),
	.w4(32'hbb97c23c),
	.w5(32'h39ae8cc2),
	.w6(32'hbbf5793f),
	.w7(32'hbc014969),
	.w8(32'h3b1697b1),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb193f2a),
	.w1(32'h3bfc8444),
	.w2(32'h3bb51aa0),
	.w3(32'hbb37e9c3),
	.w4(32'h3c02d8ac),
	.w5(32'h3c9bb5b6),
	.w6(32'h3c8bc93d),
	.w7(32'h3ca3e8fb),
	.w8(32'h3b815a05),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8468c7),
	.w1(32'hbae85801),
	.w2(32'h3c6e2f3f),
	.w3(32'h3bcce545),
	.w4(32'h3cb765ac),
	.w5(32'hba9acffc),
	.w6(32'hbc7d2a5b),
	.w7(32'h3c1087c0),
	.w8(32'hbbc16b8f),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc03d351),
	.w1(32'hbc227459),
	.w2(32'hbc7bf695),
	.w3(32'hbc3673d3),
	.w4(32'hba349da6),
	.w5(32'hbbe92184),
	.w6(32'hbc956181),
	.w7(32'hbc08c8a2),
	.w8(32'hbc0c3d05),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba7aba05),
	.w1(32'h3b2e5378),
	.w2(32'hbad865f2),
	.w3(32'h3b7822d6),
	.w4(32'h3b2890b4),
	.w5(32'hbbad3e4e),
	.w6(32'h3b9cb631),
	.w7(32'h3b67d1c4),
	.w8(32'h3bb4c406),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaaeeb88),
	.w1(32'h3b9865e1),
	.w2(32'hbb1e3cc3),
	.w3(32'hbbac6048),
	.w4(32'hbbe39934),
	.w5(32'h3b031d5e),
	.w6(32'h3b54e364),
	.w7(32'hbb577b27),
	.w8(32'h3b087463),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3fbf88),
	.w1(32'h3c39df18),
	.w2(32'h3bac30cd),
	.w3(32'hba4f4f37),
	.w4(32'h3b54e4b3),
	.w5(32'h3b53b202),
	.w6(32'hbae20229),
	.w7(32'h3ae1c4b1),
	.w8(32'hbb824656),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bad5e32),
	.w1(32'hba8aebe3),
	.w2(32'h3bc0df6b),
	.w3(32'h3ab620b4),
	.w4(32'h3bfba37c),
	.w5(32'hbc47ebc5),
	.w6(32'hbbbd149e),
	.w7(32'h3c3b35e3),
	.w8(32'hbc4574f1),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5cca4d),
	.w1(32'hbbf953d0),
	.w2(32'hbc846ba6),
	.w3(32'hbc290701),
	.w4(32'hbbe3c489),
	.w5(32'h3b8b044d),
	.w6(32'hbc8c9bf7),
	.w7(32'hbc3cd2fb),
	.w8(32'h3b6fac24),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8cce64),
	.w1(32'hbb465cb8),
	.w2(32'hbc255bbe),
	.w3(32'hbbdc54fe),
	.w4(32'h3aee67a7),
	.w5(32'h3adc4b81),
	.w6(32'hbc8e2a4f),
	.w7(32'hbb9b3cbd),
	.w8(32'hbc32c0f8),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb00d32),
	.w1(32'hbbaf8f39),
	.w2(32'h3b92d9ca),
	.w3(32'hba62c9af),
	.w4(32'h3ac72e49),
	.w5(32'hbbd01e50),
	.w6(32'hbcb60814),
	.w7(32'hba9c3711),
	.w8(32'hbbcf1f9d),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc555f83),
	.w1(32'hbc046617),
	.w2(32'hbc501c77),
	.w3(32'hbc373f7d),
	.w4(32'hbc33c4c2),
	.w5(32'hbc1f135f),
	.w6(32'hbc4a596f),
	.w7(32'hbc2d8823),
	.w8(32'hbc2f10b7),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4dd36a),
	.w1(32'hba7a1b33),
	.w2(32'hbb5e1a17),
	.w3(32'hbb17b68c),
	.w4(32'hbbec9a3a),
	.w5(32'hbbcd0570),
	.w6(32'h3b2e3280),
	.w7(32'hbaca958e),
	.w8(32'hbc15915c),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba617f1),
	.w1(32'hbc1b05d1),
	.w2(32'hb86db914),
	.w3(32'hbb6c61ab),
	.w4(32'hbb41fe09),
	.w5(32'h3b729487),
	.w6(32'hbc45819a),
	.w7(32'h3a76dfc3),
	.w8(32'h3c280655),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b274c04),
	.w1(32'h3ad2fccd),
	.w2(32'h3b2667b9),
	.w3(32'h3b956fed),
	.w4(32'h3bd8b6ba),
	.w5(32'hb9740690),
	.w6(32'hbac9f8ce),
	.w7(32'h3ae9ffb3),
	.w8(32'hbab7b69a),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb917f33),
	.w1(32'hbaf1d78b),
	.w2(32'hbb9dffeb),
	.w3(32'hba70104a),
	.w4(32'h3a4ab438),
	.w5(32'h3ae23409),
	.w6(32'h3aba1e3f),
	.w7(32'hba52f42a),
	.w8(32'h3ab950e9),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc84372d),
	.w1(32'hbb3ddef8),
	.w2(32'hbc230cfb),
	.w3(32'hbc38bb23),
	.w4(32'hba328501),
	.w5(32'hbbb95adc),
	.w6(32'hbc503f83),
	.w7(32'hbb01fa70),
	.w8(32'hbc1e8415),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc273ca4),
	.w1(32'hba93166b),
	.w2(32'hbc81b950),
	.w3(32'hbb95fcea),
	.w4(32'hbaba3879),
	.w5(32'hba980048),
	.w6(32'hbbd5c183),
	.w7(32'h38d9bfd7),
	.w8(32'hbb3b7eed),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb68444f),
	.w1(32'h3bebd0cb),
	.w2(32'hbafca85f),
	.w3(32'hbc05306a),
	.w4(32'h3b09bf2c),
	.w5(32'h3b3a5cb2),
	.w6(32'hbc8c06ef),
	.w7(32'hbb35c6d1),
	.w8(32'hbc07adf2),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4902c5),
	.w1(32'hbb982482),
	.w2(32'hbbc25055),
	.w3(32'hbb8e0b0e),
	.w4(32'hbbe0ddf9),
	.w5(32'hbabfdfde),
	.w6(32'hbc271698),
	.w7(32'hbc1d455b),
	.w8(32'h3af56a11),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39de3ef1),
	.w1(32'h3bbc85fe),
	.w2(32'hbbee4b28),
	.w3(32'h3bac2a68),
	.w4(32'hbbe4e273),
	.w5(32'h3cd6a357),
	.w6(32'h3c4ac464),
	.w7(32'hbbc43720),
	.w8(32'h3c1661e5),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb99170),
	.w1(32'hbc0babd8),
	.w2(32'h3c9e156e),
	.w3(32'hbc18e3d7),
	.w4(32'h3cc6bc1d),
	.w5(32'hbb8ef083),
	.w6(32'hbd2a63d7),
	.w7(32'h3912d11f),
	.w8(32'hba337a59),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a46684d),
	.w1(32'h3b89493e),
	.w2(32'hbbbdedd7),
	.w3(32'hbb65c9c3),
	.w4(32'hbb934bee),
	.w5(32'h3acd1965),
	.w6(32'hbc11f869),
	.w7(32'hbbf1e6cf),
	.w8(32'h3b732462),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb91cc64),
	.w1(32'h3b39e46d),
	.w2(32'hbbb37ccf),
	.w3(32'hbb649ec6),
	.w4(32'h3b45380b),
	.w5(32'h3abfc04c),
	.w6(32'hbb37e1c0),
	.w7(32'h3bf52021),
	.w8(32'hb9a61c1b),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb89c7955),
	.w1(32'hbbe902f3),
	.w2(32'hbc08899f),
	.w3(32'h3b6486ff),
	.w4(32'h3b6a8463),
	.w5(32'h3b24815c),
	.w6(32'hbc282c33),
	.w7(32'hbbe3c614),
	.w8(32'hbc0bf4e7),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9613fe),
	.w1(32'hba9cad74),
	.w2(32'hbb034510),
	.w3(32'h3b737a05),
	.w4(32'hbb886c8f),
	.w5(32'hbb858048),
	.w6(32'h3a2aca62),
	.w7(32'h38f9104d),
	.w8(32'hbc43a7fa),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3909c1),
	.w1(32'h3c1d2196),
	.w2(32'hbbcdce89),
	.w3(32'hbbb74ee9),
	.w4(32'hbc03badd),
	.w5(32'hbc1a60de),
	.w6(32'h3ba437a1),
	.w7(32'hb9ce159e),
	.w8(32'hbbcd463c),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0ac91e),
	.w1(32'hbbcbc68d),
	.w2(32'hbaf5eae6),
	.w3(32'hbc3564b5),
	.w4(32'h3b1bc7fe),
	.w5(32'hbb2d0a60),
	.w6(32'hbc805438),
	.w7(32'h3aa9e89a),
	.w8(32'hbb4daf88),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acc1215),
	.w1(32'hb7b52364),
	.w2(32'hba27d343),
	.w3(32'hbb9f4869),
	.w4(32'hba15044b),
	.w5(32'h3ac22a7d),
	.w6(32'hbc1785a5),
	.w7(32'hbba5afd9),
	.w8(32'h3a9f83ac),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b82e77d),
	.w1(32'hbabb7fbb),
	.w2(32'h3ad54f1e),
	.w3(32'hb9c458fd),
	.w4(32'hbb98777f),
	.w5(32'hbc00049f),
	.w6(32'hba776733),
	.w7(32'hba42f132),
	.w8(32'h3ae39224),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba46b64),
	.w1(32'h3bbae644),
	.w2(32'hbb5c8876),
	.w3(32'hbb0f2931),
	.w4(32'h3bd0d494),
	.w5(32'h3bbf38f1),
	.w6(32'hba890801),
	.w7(32'h3b9efffa),
	.w8(32'hbbc6f0c8),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc5d311b),
	.w1(32'h3c0272da),
	.w2(32'h3c107009),
	.w3(32'hbbeb176f),
	.w4(32'h3c620301),
	.w5(32'h3c220a8c),
	.w6(32'hbc99c2a5),
	.w7(32'h3adc5445),
	.w8(32'h3b8d2bd2),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb025d27),
	.w1(32'h3c27ee13),
	.w2(32'h3bcc35a0),
	.w3(32'hbb630b8a),
	.w4(32'h3c759a7e),
	.w5(32'hbad2f2e3),
	.w6(32'hbcd765fe),
	.w7(32'h3b6c453a),
	.w8(32'h3a0c2fae),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1b489d),
	.w1(32'hbc037cab),
	.w2(32'hba4341fc),
	.w3(32'hbc5b06da),
	.w4(32'hbb3bf4ff),
	.w5(32'h3b336dbc),
	.w6(32'hbc037e7d),
	.w7(32'hbada337b),
	.w8(32'h3a7553d2),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b888baa),
	.w1(32'h3b7f9943),
	.w2(32'h3b6b05bd),
	.w3(32'h3b5c538f),
	.w4(32'h3aa02ad9),
	.w5(32'hbb33da9a),
	.w6(32'hbac7bd5e),
	.w7(32'hba950936),
	.w8(32'hba51bb9d),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba13f507),
	.w1(32'hba87f17c),
	.w2(32'hbc035e28),
	.w3(32'hbb0fff5d),
	.w4(32'hbbca67d1),
	.w5(32'h3b8d910d),
	.w6(32'h3b865768),
	.w7(32'hbb8df87a),
	.w8(32'h3a0075f8),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c4d3e25),
	.w1(32'h3c511b5f),
	.w2(32'h3c117582),
	.w3(32'h3b972b53),
	.w4(32'h3c459a9c),
	.w5(32'hbbcb12e7),
	.w6(32'h3bd0637b),
	.w7(32'h3c06900b),
	.w8(32'hbb50e685),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2d179e),
	.w1(32'hbc00d35f),
	.w2(32'hbcb73ef9),
	.w3(32'hbbed857c),
	.w4(32'hbc61681d),
	.w5(32'hbc8757da),
	.w6(32'hbc2ac15e),
	.w7(32'hbc1f9c8b),
	.w8(32'hbc2dbf05),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf4aa76),
	.w1(32'h3c686fcf),
	.w2(32'hbc182ae5),
	.w3(32'h3bd15140),
	.w4(32'h3c03f421),
	.w5(32'h3bbfe35a),
	.w6(32'h3c9b58a3),
	.w7(32'h3c4d761e),
	.w8(32'hbb9cf9b6),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb907c2ea),
	.w1(32'h3b2283b7),
	.w2(32'h3accb923),
	.w3(32'hbb37520a),
	.w4(32'h3c4693e7),
	.w5(32'hbc0bbc3d),
	.w6(32'hbccf8536),
	.w7(32'hbb5298c3),
	.w8(32'h3a40e368),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb31fffc),
	.w1(32'h3c461f16),
	.w2(32'hbbd679ea),
	.w3(32'hb994c609),
	.w4(32'hbad245b1),
	.w5(32'h3ca464fb),
	.w6(32'h3c238388),
	.w7(32'h3b15f457),
	.w8(32'h3c00e8db),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c100eb0),
	.w1(32'hbac90fe5),
	.w2(32'hb995b6eb),
	.w3(32'h3b1d3d55),
	.w4(32'h3b7f8081),
	.w5(32'hbb570d7c),
	.w6(32'hbb0368c6),
	.w7(32'hbaf3bfa5),
	.w8(32'hbc528225),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c5c5c2f),
	.w1(32'h3bf60921),
	.w2(32'h3bd574c0),
	.w3(32'h3be98f3a),
	.w4(32'h3c424571),
	.w5(32'h3b89e466),
	.w6(32'hbba76220),
	.w7(32'h3a8968fe),
	.w8(32'h3a223218),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2f74ce),
	.w1(32'hbb5d5711),
	.w2(32'h3a98288c),
	.w3(32'hb933e3a6),
	.w4(32'h3be3631b),
	.w5(32'h3bc8af0b),
	.w6(32'hbbaeb1cf),
	.w7(32'h3b960c02),
	.w8(32'h3ab8b6be),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b341bb4),
	.w1(32'hbc399e83),
	.w2(32'h3a15a612),
	.w3(32'hbb5ebb34),
	.w4(32'hba5f3e02),
	.w5(32'hbbf3372c),
	.w6(32'hbc012f12),
	.w7(32'hbbc5026a),
	.w8(32'hbb6e9334),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd8c9b9),
	.w1(32'h3a625962),
	.w2(32'hbc2ae653),
	.w3(32'hbbc19f78),
	.w4(32'hbc318d78),
	.w5(32'hbb94061c),
	.w6(32'h39dba86d),
	.w7(32'hbbd977f3),
	.w8(32'hbaaa06b1),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe2a077),
	.w1(32'hb97c431d),
	.w2(32'hbc63bdaf),
	.w3(32'hba4042ca),
	.w4(32'hbc0de054),
	.w5(32'hbb2eb17c),
	.w6(32'h3abe2a3a),
	.w7(32'hbb9d17b6),
	.w8(32'h3b7c95ee),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc446939),
	.w1(32'h3b8388d9),
	.w2(32'hbc742033),
	.w3(32'hbb43a217),
	.w4(32'hbc15c487),
	.w5(32'hbbdd54a0),
	.w6(32'hbad897cc),
	.w7(32'hbc229d7e),
	.w8(32'hbbf5f176),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae0dc00),
	.w1(32'hbb82d0d4),
	.w2(32'hbbd2ae45),
	.w3(32'h3a02f289),
	.w4(32'hbb9341c9),
	.w5(32'hbb0e9fd3),
	.w6(32'hbbc6faae),
	.w7(32'h3abf371b),
	.w8(32'hbb5a029e),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf7ffff),
	.w1(32'hba2af28b),
	.w2(32'hb9db13c7),
	.w3(32'h3b0d80c0),
	.w4(32'h3bab9c5f),
	.w5(32'h3acbe2fc),
	.w6(32'hbc4b4152),
	.w7(32'hb90cbf00),
	.w8(32'h3a462861),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c04b54b),
	.w1(32'hba9274de),
	.w2(32'h3b982e90),
	.w3(32'h3a07dd1a),
	.w4(32'h3b8cf40b),
	.w5(32'hbac9da29),
	.w6(32'hbb9c9b3a),
	.w7(32'h3acc9d6b),
	.w8(32'h3b68ea2b),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3adae378),
	.w1(32'h3b4484a9),
	.w2(32'hbb6f5659),
	.w3(32'hb9811a41),
	.w4(32'hb9b3ee4c),
	.w5(32'h3bee10ae),
	.w6(32'hbb16b71c),
	.w7(32'hbb30f899),
	.w8(32'h3ad891fe),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b54936b),
	.w1(32'hbbd19529),
	.w2(32'hb9b0f182),
	.w3(32'hb9f89184),
	.w4(32'h3bc4404b),
	.w5(32'h3b8c2657),
	.w6(32'hbc06c3b3),
	.w7(32'h3a126039),
	.w8(32'h3b64de06),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4d7d5f),
	.w1(32'h3c6cd95a),
	.w2(32'h3c26bb4c),
	.w3(32'h3c21f81c),
	.w4(32'h3b444939),
	.w5(32'h3bcb4584),
	.w6(32'h3c99dfd1),
	.w7(32'h3bc6a136),
	.w8(32'h393463a9),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba2d126b),
	.w1(32'hbbbe3c4f),
	.w2(32'hbb5088e0),
	.w3(32'h39b3d3c6),
	.w4(32'h3c04acf9),
	.w5(32'h3a9b0b0d),
	.w6(32'hbca3e39c),
	.w7(32'hb8d32d18),
	.w8(32'hbbbeb57e),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h398780aa),
	.w1(32'hbb923ccd),
	.w2(32'hbab5d7be),
	.w3(32'hbb8848c3),
	.w4(32'h3bdba6f2),
	.w5(32'h3a20766f),
	.w6(32'hbcbfbf39),
	.w7(32'hbb8553de),
	.w8(32'hb905d3ae),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcd9318),
	.w1(32'h3bd3f77f),
	.w2(32'h3b1940bd),
	.w3(32'hb9f57d6f),
	.w4(32'hbb294802),
	.w5(32'hb999c444),
	.w6(32'hbbba7efe),
	.w7(32'h39ce87dc),
	.w8(32'h3a6b1df9),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5ed82d),
	.w1(32'hbac84fe5),
	.w2(32'hba4a2748),
	.w3(32'hbb6838da),
	.w4(32'hbb4356ab),
	.w5(32'h3b55df0e),
	.w6(32'hbc072ca7),
	.w7(32'hbb18f16a),
	.w8(32'hba5402f9),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba037d9c),
	.w1(32'hba213b4c),
	.w2(32'hbb52f7ee),
	.w3(32'h3bbb7e5b),
	.w4(32'h3b3f3df6),
	.w5(32'h389a8490),
	.w6(32'hbb1ee6c5),
	.w7(32'h3acf2ac3),
	.w8(32'h3b57f0a2),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h391a92a5),
	.w1(32'hba927bc8),
	.w2(32'hbbac3939),
	.w3(32'h39fee695),
	.w4(32'hba8a78d0),
	.w5(32'h3bb352a6),
	.w6(32'hbac26a65),
	.w7(32'h3bb61620),
	.w8(32'h3af066c8),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h397d3f56),
	.w1(32'h3b906e0f),
	.w2(32'h3b73f215),
	.w3(32'hbb4c8f5a),
	.w4(32'h3b8dea22),
	.w5(32'hbca050d6),
	.w6(32'hbb5d5f5f),
	.w7(32'h3c1e68bc),
	.w8(32'hbcbf43ec),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcb5824e),
	.w1(32'hbc8c7e32),
	.w2(32'hbd18e5df),
	.w3(32'hbc958764),
	.w4(32'hbcc36903),
	.w5(32'h398196e3),
	.w6(32'hbcb3400b),
	.w7(32'hbd06957c),
	.w8(32'hbbeb5eb8),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9c352a),
	.w1(32'h3a290924),
	.w2(32'hb8272412),
	.w3(32'hbb80ae07),
	.w4(32'h3bbb062f),
	.w5(32'hb9d2c460),
	.w6(32'hbbebe091),
	.w7(32'h3c13d8b4),
	.w8(32'h3ae3c0b3),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2e7811),
	.w1(32'h3c2258a0),
	.w2(32'hbb976447),
	.w3(32'h37fdf8f6),
	.w4(32'h3c6e07fd),
	.w5(32'hbab463a2),
	.w6(32'h3b6d5456),
	.w7(32'h3c4a5496),
	.w8(32'hbb32ca9f),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba9eb4c),
	.w1(32'h3c0914b2),
	.w2(32'h3bb584cc),
	.w3(32'hba2c7fea),
	.w4(32'hbb64f2c8),
	.w5(32'hbb262b1f),
	.w6(32'h3c663992),
	.w7(32'h3b784666),
	.w8(32'h3a31da6a),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc38378),
	.w1(32'hbb6266ac),
	.w2(32'hbb5e371a),
	.w3(32'hbba8e013),
	.w4(32'hbb887512),
	.w5(32'h3bbe32e7),
	.w6(32'hbb929bdf),
	.w7(32'h3b2e3d6a),
	.w8(32'h3a113f70),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b63422a),
	.w1(32'h3b887e69),
	.w2(32'h3c2b7a4e),
	.w3(32'h394e2e7e),
	.w4(32'h3b997b46),
	.w5(32'hbb3c749a),
	.w6(32'hbc1d2b62),
	.w7(32'h3b0a2a02),
	.w8(32'h3bc68bc6),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3ceb2e),
	.w1(32'h3b475688),
	.w2(32'hbbc05f30),
	.w3(32'hbbecd722),
	.w4(32'h3b7d4aa0),
	.w5(32'h3b45a894),
	.w6(32'hbc14023a),
	.w7(32'hbbffb0ad),
	.w8(32'hbbd1d78a),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ad8ff65),
	.w1(32'h3b3358f9),
	.w2(32'h3c38b9e4),
	.w3(32'hba6a5d6d),
	.w4(32'h3c021e93),
	.w5(32'h3b96375c),
	.w6(32'hbc797224),
	.w7(32'h3bbf6740),
	.w8(32'h3aeba0e7),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be04607),
	.w1(32'h3b31bc4e),
	.w2(32'h39bcaf42),
	.w3(32'h39fe08e6),
	.w4(32'hbb6bc938),
	.w5(32'h3b590fc8),
	.w6(32'hbb39f584),
	.w7(32'hbb6b2126),
	.w8(32'h3c0642ec),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3998a57b),
	.w1(32'hbb0292bd),
	.w2(32'hbb44a6e9),
	.w3(32'hba501314),
	.w4(32'hbb69d16e),
	.w5(32'hbc36a6bd),
	.w6(32'hbbb2583d),
	.w7(32'h3b35ed25),
	.w8(32'hbbd8c086),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc6d2544),
	.w1(32'hbb2ade2e),
	.w2(32'hbc16bdd6),
	.w3(32'hbc37e0cf),
	.w4(32'hbbe3a39a),
	.w5(32'hbbf46b7f),
	.w6(32'hbb8cd0dc),
	.w7(32'hbb2489e1),
	.w8(32'hbc0ddfee),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6129ec),
	.w1(32'hbb9ee2f1),
	.w2(32'hbc14c5b2),
	.w3(32'hbbd514a6),
	.w4(32'hba08682b),
	.w5(32'h3c2f5cb1),
	.w6(32'hbb2728cf),
	.w7(32'hbb50caa6),
	.w8(32'h3a9f6cbf),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c442e2e),
	.w1(32'hbb5209a4),
	.w2(32'h3bd41b9c),
	.w3(32'hbbadd603),
	.w4(32'h3c4e0ecd),
	.w5(32'h39304374),
	.w6(32'hbd003b4d),
	.w7(32'h386c9786),
	.w8(32'h3c6e1b60),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd2f5c8),
	.w1(32'h3beb42fd),
	.w2(32'hbb90cf6a),
	.w3(32'h3c0c2aa1),
	.w4(32'h3ba6b924),
	.w5(32'h3b0e3313),
	.w6(32'h3d1c4fcc),
	.w7(32'h3c947007),
	.w8(32'hba9aa310),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b47dd13),
	.w1(32'h3b1bdac0),
	.w2(32'h3a21cea5),
	.w3(32'h3b866b20),
	.w4(32'h3bdc68ab),
	.w5(32'hbba35398),
	.w6(32'hba56af3f),
	.w7(32'h3b14f44f),
	.w8(32'hbbd5f4f6),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb97628b),
	.w1(32'hbb20ce71),
	.w2(32'h3a8b1d52),
	.w3(32'hbafb9824),
	.w4(32'hb92fc110),
	.w5(32'hbc9712c7),
	.w6(32'hbbbd1831),
	.w7(32'h3a86152f),
	.w8(32'hbc3959c0),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbca046a6),
	.w1(32'hbb8da313),
	.w2(32'hbcd4d3e6),
	.w3(32'hbb1c8a9a),
	.w4(32'hbce5af32),
	.w5(32'h3c10f78f),
	.w6(32'h3c35e651),
	.w7(32'hbc968dbf),
	.w8(32'h3b259849),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac1a662),
	.w1(32'hbb984a58),
	.w2(32'h3a2464f6),
	.w3(32'h3b04d51b),
	.w4(32'h3a8d6e8e),
	.w5(32'h3bcf3abd),
	.w6(32'hbbc7e06f),
	.w7(32'hbb5fcbfc),
	.w8(32'hbabea447),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd3a3c9),
	.w1(32'h3b60e086),
	.w2(32'h3c09c88e),
	.w3(32'h3b551535),
	.w4(32'h3c353082),
	.w5(32'hbb9c0317),
	.w6(32'hbc957df2),
	.w7(32'h3b8343fc),
	.w8(32'h3b885821),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2fa813),
	.w1(32'h39437652),
	.w2(32'hbba6a62a),
	.w3(32'hbc2268c0),
	.w4(32'hbb8495a8),
	.w5(32'h3b0bbe82),
	.w6(32'hbb3740c1),
	.w7(32'hbb328bc2),
	.w8(32'h3a0a9a68),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b73d077),
	.w1(32'h3aff0e88),
	.w2(32'h3b08502c),
	.w3(32'hba224871),
	.w4(32'h3a04e38b),
	.w5(32'h3a9ad909),
	.w6(32'hbbf5cfe4),
	.w7(32'h3a9439cb),
	.w8(32'hbc050d76),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb788a98),
	.w1(32'hbc67cc19),
	.w2(32'hbbc5fe79),
	.w3(32'hbc1ebe92),
	.w4(32'h3900d2ea),
	.w5(32'hbb0f9d36),
	.w6(32'hbcf89e37),
	.w7(32'hbc0f6283),
	.w8(32'hb9948c54),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba67ad51),
	.w1(32'hbb4d8be0),
	.w2(32'hbaf24dec),
	.w3(32'hbb058171),
	.w4(32'hbb56c40c),
	.w5(32'hb9a47254),
	.w6(32'hbc121cf1),
	.w7(32'h3a6394f3),
	.w8(32'hbb66f715),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a0aaa2d),
	.w1(32'hbb3fdfd7),
	.w2(32'hbb5f60d4),
	.w3(32'hbc659630),
	.w4(32'hbb81732d),
	.w5(32'hbbd30d29),
	.w6(32'hbc8d2ed9),
	.w7(32'hbb9e0029),
	.w8(32'hbb1199d4),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8f187c),
	.w1(32'hbb78ff10),
	.w2(32'hbc595fc2),
	.w3(32'hbbf06d35),
	.w4(32'hbc0b4c88),
	.w5(32'hbb851eb2),
	.w6(32'h3b61685e),
	.w7(32'hbb16857f),
	.w8(32'hbc0ca1e5),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c8310),
	.w1(32'hbb912646),
	.w2(32'hbbabf2dc),
	.w3(32'h3ab23562),
	.w4(32'hbb662f00),
	.w5(32'hbbd0ae3c),
	.w6(32'h3ae4dc96),
	.w7(32'h3c027343),
	.w8(32'hbbf888b5),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc261dce),
	.w1(32'hbb672587),
	.w2(32'hbc5cc7c8),
	.w3(32'h39a7059d),
	.w4(32'hba4cc808),
	.w5(32'hba0e5fd2),
	.w6(32'hbb6c6a20),
	.w7(32'hbb51cc53),
	.w8(32'hbc0fc89a),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc149679),
	.w1(32'hbc3baf61),
	.w2(32'hbbd37900),
	.w3(32'hbc1f771b),
	.w4(32'hbad2cba6),
	.w5(32'h3b8a19c7),
	.w6(32'hbc68b440),
	.w7(32'hbb86d848),
	.w8(32'hbbfdf05f),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc38ee30),
	.w1(32'hbbb93d0e),
	.w2(32'hbbb55f36),
	.w3(32'hbba20157),
	.w4(32'hbabd33c8),
	.w5(32'hbc6a179f),
	.w6(32'hbc11e222),
	.w7(32'h3adf23aa),
	.w8(32'hbc5e7d1d),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc57b760),
	.w1(32'hbc4cba87),
	.w2(32'hbc849a36),
	.w3(32'hbbf2c2e1),
	.w4(32'hbc3b34ea),
	.w5(32'hbbad7582),
	.w6(32'hbc2c8fff),
	.w7(32'hbc73032a),
	.w8(32'hbc00a2f4),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2c8283),
	.w1(32'hbb4e1e02),
	.w2(32'hbb19d200),
	.w3(32'hbbdf11e9),
	.w4(32'hbbac2812),
	.w5(32'hbbec8439),
	.w6(32'hbc3d0ec1),
	.w7(32'hba9d57b5),
	.w8(32'hbc0de951),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb007fe8),
	.w1(32'hba75a26a),
	.w2(32'hbadbf2da),
	.w3(32'hbbf84be0),
	.w4(32'hba11751c),
	.w5(32'hbb6aa931),
	.w6(32'hbbadbaa7),
	.w7(32'hb9ebb36c),
	.w8(32'hbbd777b3),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbee5112),
	.w1(32'hbade1740),
	.w2(32'hbc098093),
	.w3(32'hbbd91a53),
	.w4(32'h3af86e82),
	.w5(32'h3b2fc9d9),
	.w6(32'hbc17ecbe),
	.w7(32'h3a7a89da),
	.w8(32'hbbc7626f),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1efd8d),
	.w1(32'h3c119b0b),
	.w2(32'h3b8b11a7),
	.w3(32'hbc1d9135),
	.w4(32'h3c7e768a),
	.w5(32'h3c369fa0),
	.w6(32'hbc4f115a),
	.w7(32'h3bf4439c),
	.w8(32'h3a328084),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0585d7),
	.w1(32'h3ac7b4bb),
	.w2(32'hbbd94dbd),
	.w3(32'hbbdc806b),
	.w4(32'h39f3a780),
	.w5(32'hbbd17214),
	.w6(32'hbc14205c),
	.w7(32'h3b37400c),
	.w8(32'hbc0366b0),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7a1c01),
	.w1(32'hba8b4228),
	.w2(32'hbb8e9264),
	.w3(32'hbb3ae187),
	.w4(32'h395c292b),
	.w5(32'hbada3516),
	.w6(32'hbac8f574),
	.w7(32'h3b9574f6),
	.w8(32'hbb8021a6),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb29bb0e),
	.w1(32'hbabcc14c),
	.w2(32'h3b61b0ca),
	.w3(32'h3a87fce0),
	.w4(32'h3ad50e25),
	.w5(32'hbb560e66),
	.w6(32'hb9752489),
	.w7(32'h3b35b566),
	.w8(32'hbc020654),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc41dc68),
	.w1(32'hbc2779c9),
	.w2(32'hbc2d27c2),
	.w3(32'hbbd8dfc7),
	.w4(32'hbb13947c),
	.w5(32'hbb729f16),
	.w6(32'hbbf9de7a),
	.w7(32'h3b32ae31),
	.w8(32'hbade382e),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb589a13),
	.w1(32'hbb1c4786),
	.w2(32'hbb8ee639),
	.w3(32'hbba9f845),
	.w4(32'hbbf33dbe),
	.w5(32'hbbf688e0),
	.w6(32'hbaf4fa02),
	.w7(32'hbb0b4856),
	.w8(32'hbb7e5288),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba77e15),
	.w1(32'hbb89e729),
	.w2(32'hbb510795),
	.w3(32'hbb3ad51f),
	.w4(32'hba9c5b7a),
	.w5(32'h3b80bc5b),
	.w6(32'hbb48daf9),
	.w7(32'hba5b5511),
	.w8(32'h3b50bbfe),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3babba18),
	.w1(32'h3bd8aa30),
	.w2(32'h3bd46fe4),
	.w3(32'h3bd37bff),
	.w4(32'h3bb85e59),
	.w5(32'h3a8ab431),
	.w6(32'hba9f9ad4),
	.w7(32'h3b036401),
	.w8(32'h38905780),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfe0ff0),
	.w1(32'hbc084828),
	.w2(32'hbc07b0aa),
	.w3(32'hbc09f59f),
	.w4(32'hbb93a277),
	.w5(32'hbbc17159),
	.w6(32'hbc01b10c),
	.w7(32'hbbb4894f),
	.w8(32'hbbe8dcfa),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b176d53),
	.w1(32'h3bcedc34),
	.w2(32'hbae21022),
	.w3(32'hbb091fc2),
	.w4(32'h3b7779f2),
	.w5(32'hbb8d7ecf),
	.w6(32'hbbba5191),
	.w7(32'h37202cc6),
	.w8(32'hbbd82ba4),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4e5439),
	.w1(32'h3ac70d8a),
	.w2(32'hbb28e2ea),
	.w3(32'hbc041d16),
	.w4(32'hbaebf7e7),
	.w5(32'h3ac2af21),
	.w6(32'hbbc08e88),
	.w7(32'hbb2410cd),
	.w8(32'hbb4519ce),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf6638c),
	.w1(32'hbae8cb5e),
	.w2(32'hbbe98b6e),
	.w3(32'hb9f56cf8),
	.w4(32'h3ad4d4ff),
	.w5(32'hbb345bf0),
	.w6(32'hbb38ddd4),
	.w7(32'hba30fc50),
	.w8(32'hba1c238f),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae5a15d),
	.w1(32'h3b5e7cda),
	.w2(32'h3aee7cb3),
	.w3(32'hb79a2500),
	.w4(32'h3b8543c1),
	.w5(32'hbada3f3e),
	.w6(32'hba2741c1),
	.w7(32'h3b4fa89f),
	.w8(32'hb8d352be),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd72a87),
	.w1(32'hbb81b527),
	.w2(32'hbbb8572a),
	.w3(32'hbb22a4d9),
	.w4(32'h3a4a1cb6),
	.w5(32'hbb903bf5),
	.w6(32'hbb22f205),
	.w7(32'h397a9222),
	.w8(32'hbbd1feb1),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc03c4f7),
	.w1(32'hba88688c),
	.w2(32'hbbf35fcf),
	.w3(32'hbbdd7104),
	.w4(32'hb880fbd0),
	.w5(32'hba505daa),
	.w6(32'hbb7ed56c),
	.w7(32'hbb02acb4),
	.w8(32'hbb8c1784),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb94cb202),
	.w1(32'hba86c3ce),
	.w2(32'hbb03a41a),
	.w3(32'hba94b195),
	.w4(32'hbb3b84af),
	.w5(32'h3b8e8025),
	.w6(32'hbb14aa82),
	.w7(32'hbabf92aa),
	.w8(32'h3b8209e4),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b966275),
	.w1(32'h3bd7f480),
	.w2(32'h39c85a6f),
	.w3(32'h3b902106),
	.w4(32'h3ad5781a),
	.w5(32'hbbc7076d),
	.w6(32'h3bb94ed7),
	.w7(32'h3a1b09b9),
	.w8(32'hbbb6c174),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8cfbe5),
	.w1(32'hbc1333e2),
	.w2(32'hbb3083c1),
	.w3(32'hbbdaff32),
	.w4(32'hbb82ed83),
	.w5(32'h3b1af3c0),
	.w6(32'hbbc28519),
	.w7(32'hbb5acdb5),
	.w8(32'h3b70729e),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b173eb5),
	.w1(32'h3a2e455d),
	.w2(32'h3a0f314c),
	.w3(32'hba9e6726),
	.w4(32'hb8c026df),
	.w5(32'hbb7be60d),
	.w6(32'h3a697677),
	.w7(32'h3ab68647),
	.w8(32'hbbbbc057),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe8b8e2),
	.w1(32'hbb9b212b),
	.w2(32'hbbab984e),
	.w3(32'hbc1d9888),
	.w4(32'hbb0bb6c7),
	.w5(32'h3adc181c),
	.w6(32'hbc203c5b),
	.w7(32'hbb35b9c7),
	.w8(32'hbb0fd95d),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb7daef3c),
	.w1(32'hbacc4d50),
	.w2(32'hbb46e126),
	.w3(32'h3b50e7c5),
	.w4(32'h3abe3d69),
	.w5(32'hbb7bdd68),
	.w6(32'h3b0460b7),
	.w7(32'h3a066c19),
	.w8(32'hba9fc276),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba58ad1),
	.w1(32'hbb0f5def),
	.w2(32'hbb679b89),
	.w3(32'hbb430ab6),
	.w4(32'hbb49e966),
	.w5(32'hbc10bcb6),
	.w6(32'h3bc15f69),
	.w7(32'hb9823242),
	.w8(32'hbba78a7a),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc26e63f),
	.w1(32'hbbb0c935),
	.w2(32'hbbf4ab0c),
	.w3(32'hbc3f12b4),
	.w4(32'hbb89e469),
	.w5(32'hbb4e569d),
	.w6(32'hbc5475fd),
	.w7(32'hbb8d3670),
	.w8(32'hbb0746c5),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39f5d6fd),
	.w1(32'h3a948040),
	.w2(32'hbaa3aa6a),
	.w3(32'hba7658a7),
	.w4(32'hb9c1eac0),
	.w5(32'hbb1125d8),
	.w6(32'h39d087f1),
	.w7(32'hba40bcea),
	.w8(32'hbb27cee5),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38e8408e),
	.w1(32'hbb8b95ff),
	.w2(32'hbbba5ece),
	.w3(32'hbba6bed6),
	.w4(32'hbb7978b2),
	.w5(32'h3a730071),
	.w6(32'hbbbaae49),
	.w7(32'hbb9253d3),
	.w8(32'hb9b094cd),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8cab8f),
	.w1(32'hbb904f3a),
	.w2(32'hbb3a7865),
	.w3(32'h3882cc1b),
	.w4(32'hba10851f),
	.w5(32'h3ae298b9),
	.w6(32'hb95dbb39),
	.w7(32'hba0cfcb9),
	.w8(32'hb907c00f),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3beb633a),
	.w1(32'h3be3c736),
	.w2(32'h3b48abe0),
	.w3(32'hba86b77a),
	.w4(32'hbb36b04c),
	.w5(32'h3ab1b8d5),
	.w6(32'hbbb13475),
	.w7(32'hbbb18138),
	.w8(32'hba22b326),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad95678),
	.w1(32'hbb85ba5f),
	.w2(32'hbbdca7ec),
	.w3(32'h3aac53e4),
	.w4(32'h399ce33d),
	.w5(32'hbb972571),
	.w6(32'h3a888f16),
	.w7(32'hb9b9d754),
	.w8(32'hbb7c7ee7),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4abfc1),
	.w1(32'h3b8ee90e),
	.w2(32'hbaca64ce),
	.w3(32'hbae21eea),
	.w4(32'h3aeb4403),
	.w5(32'hbc4dff2a),
	.w6(32'hba4b5f16),
	.w7(32'h3b173f5a),
	.w8(32'hbc0a8efd),
)
Conv2D3x3_Inst128(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4127:4096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst128_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba29894d),
	.w1(32'hbb9b0324),
	.w2(32'hbb966a80),
	.w3(32'hbbba89fa),
	.w4(32'hbc004f96),
	.w5(32'h3b80e2ea),
	.w6(32'hbae8005b),
	.w7(32'hbb6a9fcb),
	.w8(32'hbaf8eeb0),
)
Conv2D3x3_Inst129(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4159:4128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst129_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb16f77),
	.w1(32'h39e6e8ce),
	.w2(32'h3a80a3e2),
	.w3(32'hbb5ff147),
	.w4(32'hbae2d6bc),
	.w5(32'hbb363da3),
	.w6(32'hbb94448c),
	.w7(32'hba9f9278),
	.w8(32'hbafa3cf8),
)
Conv2D3x3_Inst130(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4191:4160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst130_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39e24513),
	.w1(32'h3b11f3f9),
	.w2(32'h3b07a4e9),
	.w3(32'hbb405d4d),
	.w4(32'h38e4fa8d),
	.w5(32'h3a2e60d4),
	.w6(32'h3a47b4fc),
	.w7(32'h3b1209d4),
	.w8(32'hbb9a9572),
)
Conv2D3x3_Inst131(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4223:4192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst131_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba38f478),
	.w1(32'hbb4cd529),
	.w2(32'hbbb01f45),
	.w3(32'hba8c050f),
	.w4(32'h3b310986),
	.w5(32'hbab43df5),
	.w6(32'hbc133324),
	.w7(32'hbbb9b376),
	.w8(32'hbb57f51d),
)
Conv2D3x3_Inst132(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4255:4224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst132_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb6a0528),
	.w1(32'h3903cd79),
	.w2(32'hbb6468ed),
	.w3(32'hbb736316),
	.w4(32'h3a56138c),
	.w5(32'hbb056f1d),
	.w6(32'hbba2477d),
	.w7(32'hba1c57e1),
	.w8(32'hbb21323a),
)
Conv2D3x3_Inst133(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4287:4256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst133_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba83f6c5),
	.w1(32'hb93fd30d),
	.w2(32'hbc1b4335),
	.w3(32'hbbc62d15),
	.w4(32'hbbc405af),
	.w5(32'hbc122e4b),
	.w6(32'hbb851ce2),
	.w7(32'hbc126221),
	.w8(32'hbc58f1a9),
)
Conv2D3x3_Inst134(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4319:4288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst134_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc97e36),
	.w1(32'h3bb79136),
	.w2(32'hbafc6e51),
	.w3(32'hbb914488),
	.w4(32'h3c08d67c),
	.w5(32'h3b0b566b),
	.w6(32'h3a261ac5),
	.w7(32'h3c037d97),
	.w8(32'h388d1f1d),
)
Conv2D3x3_Inst135(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4351:4320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst135_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9dc0ca),
	.w1(32'h3baa626f),
	.w2(32'hba845397),
	.w3(32'h3a090d31),
	.w4(32'h3b6b84bf),
	.w5(32'hba347e01),
	.w6(32'h3af87a5a),
	.w7(32'h3afea85d),
	.w8(32'hbb32f26a),
)
Conv2D3x3_Inst136(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4383:4352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst136_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac970a6),
	.w1(32'h3abd98d6),
	.w2(32'hbb908e39),
	.w3(32'hbb19bc84),
	.w4(32'hba7f0777),
	.w5(32'hbc22b9ad),
	.w6(32'hbacf505e),
	.w7(32'hbaddb958),
	.w8(32'hbc1a0fc8),
)
Conv2D3x3_Inst137(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4415:4384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst137_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbec01a0),
	.w1(32'h3a20fb37),
	.w2(32'hba9a7bed),
	.w3(32'hbb5a6e0e),
	.w4(32'h3aae859b),
	.w5(32'h388a680b),
	.w6(32'hbbc38523),
	.w7(32'hbafffc81),
	.w8(32'hbb3385b6),
)
Conv2D3x3_Inst138(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4447:4416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst138_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbfa19ef),
	.w1(32'hba8c813f),
	.w2(32'hbb736ed5),
	.w3(32'hba982f03),
	.w4(32'h3b6dc5f2),
	.w5(32'hbc1a337e),
	.w6(32'hbaf58a86),
	.w7(32'h39ccb8c6),
	.w8(32'hbc0adb3f),
)
Conv2D3x3_Inst139(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4479:4448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst139_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb827be6),
	.w1(32'hbb695fd4),
	.w2(32'hbbfdcf61),
	.w3(32'hbb8840aa),
	.w4(32'hbb8ebd02),
	.w5(32'hba3bb14d),
	.w6(32'hbbd05c2a),
	.w7(32'hbb9a36f7),
	.w8(32'hba40260a),
)
Conv2D3x3_Inst140(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4511:4480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst140_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0406fa),
	.w1(32'h3b66efe5),
	.w2(32'hbb9e1103),
	.w3(32'hbc3f18e6),
	.w4(32'h3ac029f0),
	.w5(32'hbb4da34b),
	.w6(32'hbbe01233),
	.w7(32'h39b1f794),
	.w8(32'hbbb41803),
)
Conv2D3x3_Inst141(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4543:4512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst141_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa0e5f5),
	.w1(32'h3b5c392a),
	.w2(32'h3b456851),
	.w3(32'hbb96bf1a),
	.w4(32'hbab24b83),
	.w5(32'hbb18c6c8),
	.w6(32'hbb9238a2),
	.w7(32'hba06d749),
	.w8(32'hbb201283),
)
Conv2D3x3_Inst142(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4575:4544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst142_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3acb5d07),
	.w1(32'hbaa004c9),
	.w2(32'hbb916ef8),
	.w3(32'h394aced7),
	.w4(32'hbb6f0391),
	.w5(32'h3793900e),
	.w6(32'h3b60bebf),
	.w7(32'hbb467823),
	.w8(32'h3a265b2c),
)
Conv2D3x3_Inst143(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4607:4576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst143_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba8ce46),
	.w1(32'h38a2f11f),
	.w2(32'h3b6ad982),
	.w3(32'h3a29d1f6),
	.w4(32'hbb19e5cb),
	.w5(32'hbabd54d9),
	.w6(32'hbb400b6d),
	.w7(32'hba3687a4),
	.w8(32'hb8c80d43),
)
Conv2D3x3_Inst144(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4639:4608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst144_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbadcb5a7),
	.w1(32'h3988b007),
	.w2(32'hba6234f3),
	.w3(32'hbb6c3af2),
	.w4(32'hbb2c054c),
	.w5(32'hb8a27700),
	.w6(32'hba5020dc),
	.w7(32'hba93431d),
	.w8(32'hba1dd8b6),
)
Conv2D3x3_Inst145(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4671:4640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst145_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc2364c),
	.w1(32'h38d0d2bf),
	.w2(32'hbabd2a4e),
	.w3(32'hbbec8020),
	.w4(32'h399f6a22),
	.w5(32'hbb862301),
	.w6(32'hbbb7df5a),
	.w7(32'h39429e5b),
	.w8(32'hbbcd4295),
)
Conv2D3x3_Inst146(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4703:4672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst146_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc48f48b),
	.w1(32'hbc1c82c4),
	.w2(32'hbc282761),
	.w3(32'hbc70ea11),
	.w4(32'hbbd301eb),
	.w5(32'hbc02b39b),
	.w6(32'hbc455a13),
	.w7(32'hbc0e6dae),
	.w8(32'hbbf20c3c),
)
Conv2D3x3_Inst147(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4735:4704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst147_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97c0006),
	.w1(32'h3bceed43),
	.w2(32'hba89e202),
	.w3(32'h3b955493),
	.w4(32'hbb3e84fd),
	.w5(32'h3b5d2bf4),
	.w6(32'h3c107d37),
	.w7(32'h3a8310e7),
	.w8(32'h3b73b28a),
)
Conv2D3x3_Inst148(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4767:4736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst148_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b061055),
	.w1(32'h3a739506),
	.w2(32'hbbcd2b24),
	.w3(32'hba2d749c),
	.w4(32'h3a8128ce),
	.w5(32'hbc2467f3),
	.w6(32'hbb205640),
	.w7(32'h3992ef85),
	.w8(32'hbbeb2687),
)
Conv2D3x3_Inst149(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4799:4768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst149_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbde9e9e),
	.w1(32'hbb36034a),
	.w2(32'hbb8da975),
	.w3(32'hbb962a88),
	.w4(32'hbacb5120),
	.w5(32'hbbed4cf7),
	.w6(32'hbb04dc93),
	.w7(32'hba6381af),
	.w8(32'hbc10179d),
)
Conv2D3x3_Inst150(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4831:4800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst150_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb784a2d),
	.w1(32'h3bb358e9),
	.w2(32'hbc10bf4e),
	.w3(32'hbbb4668b),
	.w4(32'hbbe1ed9b),
	.w5(32'hbbdbd044),
	.w6(32'h3be8bf20),
	.w7(32'hbb713b05),
	.w8(32'hbbab9bc2),
)
Conv2D3x3_Inst151(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4863:4832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst151_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8e4bc2),
	.w1(32'h3b9a9d7f),
	.w2(32'hbb43b6a9),
	.w3(32'hbbcc7fd8),
	.w4(32'hb916fde4),
	.w5(32'h3a01db1d),
	.w6(32'hbb976031),
	.w7(32'h3b84fda0),
	.w8(32'hbb98634d),
)
Conv2D3x3_Inst152(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4895:4864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst152_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8641cd),
	.w1(32'h3bbf4fbc),
	.w2(32'h3b86179f),
	.w3(32'h3a9b30da),
	.w4(32'h3b203282),
	.w5(32'h3b03c23a),
	.w6(32'hbb4818c9),
	.w7(32'hbab586ae),
	.w8(32'h38a9b061),
)
Conv2D3x3_Inst153(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4927:4896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst153_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae3b3fd),
	.w1(32'hba4c5c1d),
	.w2(32'hbaab3d95),
	.w3(32'hb8d6db05),
	.w4(32'hbabf7e6c),
	.w5(32'h3b87db25),
	.w6(32'hb9d2fb13),
	.w7(32'hbb101043),
	.w8(32'h3b868aa8),
)
Conv2D3x3_Inst154(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4959:4928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst154_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b9a299e),
	.w1(32'h3c1342c0),
	.w2(32'h3b33d987),
	.w3(32'h3a91d171),
	.w4(32'h3bf42dd5),
	.w5(32'hba99c819),
	.w6(32'hbb800c29),
	.w7(32'h3b234a27),
	.w8(32'h3a8dde64),
)
Conv2D3x3_Inst155(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4991:4960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst155_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbcecbf5),
	.w1(32'h3b3de66f),
	.w2(32'h3a00ea93),
	.w3(32'hbc2e0675),
	.w4(32'hba84c4da),
	.w5(32'h3ac8bbe7),
	.w6(32'hbbecfab5),
	.w7(32'hba54ea29),
	.w8(32'hbab3f9ea),
)
Conv2D3x3_Inst156(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5023:4992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst156_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaf1a17a),
	.w1(32'h3b887f1a),
	.w2(32'h3a0b2995),
	.w3(32'hbb4722fc),
	.w4(32'h3b0b7dd2),
	.w5(32'hbb7588f8),
	.w6(32'hbae4a5ef),
	.w7(32'h3b6b5549),
	.w8(32'hbc0a8d11),
)
Conv2D3x3_Inst157(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5055:5024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst157_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb394b46),
	.w1(32'hbae2a2ec),
	.w2(32'hbc09814c),
	.w3(32'hbbbb5d3c),
	.w4(32'hbbbe65c6),
	.w5(32'h395c0d1b),
	.w6(32'hbba22cec),
	.w7(32'hbc0a9134),
	.w8(32'h3acd5da7),
)
Conv2D3x3_Inst158(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5087:5056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst158_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb54536a),
	.w1(32'h3af3b054),
	.w2(32'hbb4e30cd),
	.w3(32'h3b069f37),
	.w4(32'h3b0cbb3a),
	.w5(32'h3b3be8a5),
	.w6(32'h3b676a0f),
	.w7(32'h3ae0b790),
	.w8(32'hbac84416),
)
Conv2D3x3_Inst159(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5119:5088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst159_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3488bd),
	.w1(32'hbb7cc3ae),
	.w2(32'hbadb5ef1),
	.w3(32'hbb849712),
	.w4(32'hba079b24),
	.w5(32'hbbbe5a24),
	.w6(32'hbb9855f1),
	.w7(32'h3a0fdaa1),
	.w8(32'hbb9fb27d),
)
Conv2D3x3_Inst160(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5151:5120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst160_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba91392f),
	.w1(32'hba611504),
	.w2(32'hbae8d19f),
	.w3(32'hbabeb8c3),
	.w4(32'hbb5a759d),
	.w5(32'hbb8019da),
	.w6(32'hba9863d1),
	.w7(32'hbad16f36),
	.w8(32'hbafa1bb5),
)
Conv2D3x3_Inst161(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5183:5152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst161_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb869bbb),
	.w1(32'hba0e2543),
	.w2(32'hbb23b181),
	.w3(32'hbafbcb08),
	.w4(32'h3b70b5f3),
	.w5(32'hbb5549be),
	.w6(32'hba9d172b),
	.w7(32'h3b347f5c),
	.w8(32'hbbac5b42),
)
Conv2D3x3_Inst162(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5215:5184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst162_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2361de),
	.w1(32'h3b07b329),
	.w2(32'hb8171dde),
	.w3(32'hbb84d5f3),
	.w4(32'hbb2e95e8),
	.w5(32'hbb2a8f1c),
	.w6(32'hbace1ec8),
	.w7(32'hba11cec7),
	.w8(32'hbbae8e9c),
)
Conv2D3x3_Inst163(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5247:5216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst163_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad4c9d3),
	.w1(32'hbc1225f8),
	.w2(32'hbbe05012),
	.w3(32'hbb3b2214),
	.w4(32'hbb9ea74e),
	.w5(32'hbbb6bef3),
	.w6(32'hbbc265e1),
	.w7(32'hbbf9ffde),
	.w8(32'hbbe5bfa0),
)
Conv2D3x3_Inst164(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5279:5248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst164_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba878fe1),
	.w1(32'h3a70888d),
	.w2(32'hbb5f9a41),
	.w3(32'hbaa49eb2),
	.w4(32'hbb1f6e05),
	.w5(32'hbbaaa1a5),
	.w6(32'h3b940bb6),
	.w7(32'hbb532066),
	.w8(32'hbb2ce1eb),
)
Conv2D3x3_Inst165(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5311:5280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst165_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aadea0e),
	.w1(32'h3a820794),
	.w2(32'h3b264f14),
	.w3(32'hbbb0d4a4),
	.w4(32'hbad79452),
	.w5(32'h3b8deda2),
	.w6(32'hbb7e8195),
	.w7(32'hbaa519a8),
	.w8(32'h3b0c3683),
)
Conv2D3x3_Inst166(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5343:5312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst166_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb967694),
	.w1(32'hbb2c47b7),
	.w2(32'hbadedcf9),
	.w3(32'h3bc08fcb),
	.w4(32'h3bb71c53),
	.w5(32'h39cd8dee),
	.w6(32'h3b293e13),
	.w7(32'h3b76a2e2),
	.w8(32'hb810be1e),
)
Conv2D3x3_Inst167(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5375:5344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst167_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc85246),
	.w1(32'hbb4ca346),
	.w2(32'hbbf873e5),
	.w3(32'hbb685015),
	.w4(32'h3a66ae38),
	.w5(32'hbbba0ad4),
	.w6(32'hbb795e55),
	.w7(32'h3ab332ef),
	.w8(32'hbbe5f2f1),
)
Conv2D3x3_Inst168(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5407:5376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst168_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c193c05),
	.w1(32'h3c282fa4),
	.w2(32'h3bc3614a),
	.w3(32'h3bb76e25),
	.w4(32'h3b88881a),
	.w5(32'hbb2f3a0d),
	.w6(32'h3ac67bbe),
	.w7(32'h3978f5a8),
	.w8(32'hb9d9650b),
)
Conv2D3x3_Inst169(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5439:5408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst169_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd5c059),
	.w1(32'hbadac7a0),
	.w2(32'hbbf5c955),
	.w3(32'hbbac5851),
	.w4(32'hb89c2cf4),
	.w5(32'hbc2593c6),
	.w6(32'h3b1e2fcc),
	.w7(32'h3a2520a6),
	.w8(32'hbc611635),
)
Conv2D3x3_Inst170(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5471:5440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst170_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc1fa37b),
	.w1(32'hbc26e62d),
	.w2(32'hbc03f096),
	.w3(32'hbc3ddaef),
	.w4(32'hbbdc11d8),
	.w5(32'hbb151a36),
	.w6(32'hbc392463),
	.w7(32'hbc0dd5c2),
	.w8(32'hbb86180a),
)
Conv2D3x3_Inst171(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5503:5472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst171_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc108b41),
	.w1(32'hbad59246),
	.w2(32'hbbbbc65f),
	.w3(32'hbc57c8b5),
	.w4(32'hbb6bb3a7),
	.w5(32'hbc0b6a66),
	.w6(32'hbc493371),
	.w7(32'hbbb1b42a),
	.w8(32'hbc827576),
)
Conv2D3x3_Inst172(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5535:5504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst172_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b22fe9b),
	.w1(32'h3bb327c5),
	.w2(32'h3b260700),
	.w3(32'hbc20293b),
	.w4(32'hba9506a9),
	.w5(32'hbb7afec4),
	.w6(32'hbcbc8b98),
	.w7(32'hbbb4119d),
	.w8(32'hbbd400b4),
)
Conv2D3x3_Inst173(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5567:5536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst173_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb916ca9),
	.w1(32'hbbeaded7),
	.w2(32'hbc250cdd),
	.w3(32'hbbb23093),
	.w4(32'hbb85c93e),
	.w5(32'hbb79ccdf),
	.w6(32'hbc16bc58),
	.w7(32'hbbb25f1f),
	.w8(32'h3a09ebd5),
)
Conv2D3x3_Inst174(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5599:5568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst174_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf7d5c1),
	.w1(32'h3bc59c1a),
	.w2(32'h3ba60e8f),
	.w3(32'h3bb42498),
	.w4(32'h3b3fdfb6),
	.w5(32'hbbb478fe),
	.w6(32'h3bf97746),
	.w7(32'h3ba21723),
	.w8(32'hbbc04c26),
)
Conv2D3x3_Inst175(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5631:5600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst175_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb45bb86),
	.w1(32'h3b08c99e),
	.w2(32'hbbab6f60),
	.w3(32'hbb91df2e),
	.w4(32'hbb29d8d6),
	.w5(32'h3b704540),
	.w6(32'hbaa1cbde),
	.w7(32'hbb8e8068),
	.w8(32'h3b5c25e4),
)
Conv2D3x3_Inst176(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5663:5632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst176_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf6cc84),
	.w1(32'h3b61c3eb),
	.w2(32'h3a2af5cb),
	.w3(32'h3b3ff39a),
	.w4(32'h3a716ce1),
	.w5(32'h3aab491c),
	.w6(32'h3b44b8ec),
	.w7(32'hb9e8438a),
	.w8(32'hbad88e47),
)
Conv2D3x3_Inst177(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5695:5664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst177_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb2040cb),
	.w1(32'hbbd693be),
	.w2(32'hbb9ce7f7),
	.w3(32'hba47616f),
	.w4(32'hba9ef997),
	.w5(32'hbb815879),
	.w6(32'hbb5e9ff4),
	.w7(32'hbb3d20b1),
	.w8(32'hbb1825b5),
)
Conv2D3x3_Inst178(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5727:5696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst178_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb66ec6f),
	.w1(32'hbb34bc42),
	.w2(32'hba4b27a4),
	.w3(32'hbb4de4fb),
	.w4(32'hb81cc231),
	.w5(32'h3a02fc63),
	.w6(32'hba4140c9),
	.w7(32'hb8e47b4f),
	.w8(32'hbb95787d),
)
Conv2D3x3_Inst179(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5759:5728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst179_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc232cc9),
	.w1(32'hbbd624ce),
	.w2(32'hbc2cb98b),
	.w3(32'hbb8ebdfb),
	.w4(32'hbb06e3c5),
	.w5(32'hbb8e057b),
	.w6(32'hbbd053d2),
	.w7(32'hbbe38a77),
	.w8(32'hbb9de72c),
)
Conv2D3x3_Inst180(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5791:5760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst180_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb00d99b),
	.w1(32'hbb9241fc),
	.w2(32'h3b398b65),
	.w3(32'hbac1c640),
	.w4(32'h38b42cfe),
	.w5(32'hb97f6c7d),
	.w6(32'hbb1f76e4),
	.w7(32'hbaf11d2e),
	.w8(32'hba8098be),
)
Conv2D3x3_Inst181(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5823:5792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst181_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a5cc9d7),
	.w1(32'h3994f534),
	.w2(32'hba02b9f8),
	.w3(32'h3a9d1a54),
	.w4(32'h3aeb5e41),
	.w5(32'hbb240f7b),
	.w6(32'hbaccb256),
	.w7(32'hbae4390e),
	.w8(32'hba48df58),
)
Conv2D3x3_Inst182(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5855:5824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst182_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb62cac4),
	.w1(32'hb9808691),
	.w2(32'hbb273c22),
	.w3(32'hbb610613),
	.w4(32'hbaa32134),
	.w5(32'h3b30b8a4),
	.w6(32'hba98783c),
	.w7(32'hbacbe275),
	.w8(32'h3b3edb58),
)
Conv2D3x3_Inst183(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5887:5856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst183_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9eb7677),
	.w1(32'h3b0423cd),
	.w2(32'hba78b55a),
	.w3(32'hba494079),
	.w4(32'h3b9d2229),
	.w5(32'hbb4c7fde),
	.w6(32'hbabd5e91),
	.w7(32'h3b38cff4),
	.w8(32'hbba5f17e),
)
Conv2D3x3_Inst184(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5919:5888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst184_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3141dc),
	.w1(32'hbb11792b),
	.w2(32'hbb2ec43f),
	.w3(32'hbaa5e44b),
	.w4(32'h3b44b849),
	.w5(32'h3b9564dc),
	.w6(32'hb8c0ce66),
	.w7(32'h3bb6f363),
	.w8(32'h3b95398e),
)
Conv2D3x3_Inst185(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5951:5920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst185_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb6f2c8),
	.w1(32'h3bb5ba98),
	.w2(32'hb827c56e),
	.w3(32'h3b891e65),
	.w4(32'h3b021e2b),
	.w5(32'h3bcb89a3),
	.w6(32'h3bd68a9e),
	.w7(32'hbae95a89),
	.w8(32'h3a768fda),
)
Conv2D3x3_Inst186(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[5983:5952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst186_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb959d319),
	.w1(32'hbc0e212e),
	.w2(32'hbc47ae99),
	.w3(32'h3a8ac608),
	.w4(32'h3adc61f6),
	.w5(32'hbc0608f9),
	.w6(32'hbbff778c),
	.w7(32'hba4ea49c),
	.w8(32'hbb81b0d6),
)
Conv2D3x3_Inst187(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6015:5984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst187_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdafad5),
	.w1(32'h3b5c8e26),
	.w2(32'hbba72214),
	.w3(32'hbc25a963),
	.w4(32'h3baa0d36),
	.w5(32'hba11b343),
	.w6(32'hbbfad860),
	.w7(32'h3a5976d5),
	.w8(32'hbbd2b466),
)
Conv2D3x3_Inst188(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6047:6016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst188_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6caef2),
	.w1(32'hbad0f914),
	.w2(32'hbb3c4aa7),
	.w3(32'hbb46bf03),
	.w4(32'hbb6bc445),
	.w5(32'hbb215b29),
	.w6(32'hbbff6804),
	.w7(32'hbbf82ee8),
	.w8(32'hbb7addc2),
)
Conv2D3x3_Inst189(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6079:6048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst189_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba717c35),
	.w1(32'hbaca523c),
	.w2(32'hbadbbc9f),
	.w3(32'h3a344287),
	.w4(32'h3b0f18b8),
	.w5(32'hbaa245c3),
	.w6(32'hbb2381be),
	.w7(32'hbb24e023),
	.w8(32'hba0002e8),
)
Conv2D3x3_Inst190(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6111:6080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst190_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb014307),
	.w1(32'h39b3c866),
	.w2(32'h39a54473),
	.w3(32'hba566b5c),
	.w4(32'h3a130024),
	.w5(32'hbb377b39),
	.w6(32'h3aa17dd5),
	.w7(32'hb929f0e1),
	.w8(32'hbb8f19b9),
)
Conv2D3x3_Inst191(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6143:6112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst191_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb718e92),
	.w1(32'hbaf58e54),
	.w2(32'h3ac5ac49),
	.w3(32'hbb4c9db6),
	.w4(32'h3ae5fceb),
	.w5(32'hba99c911),
	.w6(32'hbb5665ea),
	.w7(32'hba9cd373),
	.w8(32'hba8031d4),
)
Conv2D3x3_Inst192(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6175:6144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst192_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba24d43f),
	.w1(32'hbb783966),
	.w2(32'hbbaf4ec7),
	.w3(32'h3aa35b0d),
	.w4(32'h3ae520e0),
	.w5(32'hbb869882),
	.w6(32'hbb35bc1a),
	.w7(32'hbb62ea16),
	.w8(32'hbbb1aa3a),
)
Conv2D3x3_Inst193(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6207:6176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst193_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb1e039),
	.w1(32'h3b75f389),
	.w2(32'hba35fe51),
	.w3(32'hbaabf274),
	.w4(32'h3b63b331),
	.w5(32'hbb8eea6a),
	.w6(32'hbb8ba29b),
	.w7(32'h3b34c281),
	.w8(32'hbc15c98b),
)
Conv2D3x3_Inst194(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6239:6208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst194_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbf3da0d),
	.w1(32'h3b802238),
	.w2(32'h3af55713),
	.w3(32'hbb9e346f),
	.w4(32'h3b92fb3c),
	.w5(32'h38095dce),
	.w6(32'hbbf767e1),
	.w7(32'h3b3f1427),
	.w8(32'hbbb5a6bf),
)
Conv2D3x3_Inst195(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6271:6240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst195_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1e8600),
	.w1(32'hb9f383cb),
	.w2(32'hb9ed81fa),
	.w3(32'hbb77122f),
	.w4(32'h3aa4e980),
	.w5(32'h39d5d7da),
	.w6(32'hbb28ff27),
	.w7(32'h39520bd5),
	.w8(32'hbb0f7f20),
)
Conv2D3x3_Inst196(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6303:6272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst196_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb1f6a0),
	.w1(32'hbb87c6e1),
	.w2(32'hbc307017),
	.w3(32'hbc14cc8c),
	.w4(32'hbb51aa7b),
	.w5(32'hbbdad2bb),
	.w6(32'hbc0621a5),
	.w7(32'hbb8c75ce),
	.w8(32'hbc27709f),
)
Conv2D3x3_Inst197(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6335:6304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst197_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaae828c),
	.w1(32'hbb1c5be1),
	.w2(32'hbb0e9089),
	.w3(32'hbb8ee5c1),
	.w4(32'hbb9483e7),
	.w5(32'hbbac5fc0),
	.w6(32'hbb286b35),
	.w7(32'hbb9c3e9b),
	.w8(32'hbbd93899),
)
Conv2D3x3_Inst198(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6367:6336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst198_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb45e3b7),
	.w1(32'h3bc1ca98),
	.w2(32'hb947d068),
	.w3(32'h3a030281),
	.w4(32'hb9608b44),
	.w5(32'hbb84dcda),
	.w6(32'h3b754f2e),
	.w7(32'h3b1ca8b5),
	.w8(32'hbb0d94bb),
)
Conv2D3x3_Inst199(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6399:6368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst199_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4f5adb),
	.w1(32'h3acd1c99),
	.w2(32'h3ba1e8a5),
	.w3(32'hbbe7bcf8),
	.w4(32'hba7f3000),
	.w5(32'hbb5e387a),
	.w6(32'hbaff30e9),
	.w7(32'h3adee6d0),
	.w8(32'hba4c8884),
)
Conv2D3x3_Inst200(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6431:6400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst200_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb093681),
	.w1(32'hbb2cc3e7),
	.w2(32'h3a17d306),
	.w3(32'hbb94bd05),
	.w4(32'hbb6fc595),
	.w5(32'hbb4b6411),
	.w6(32'hbb2cf7d4),
	.w7(32'hbb239a39),
	.w8(32'hba2256a7),
)
Conv2D3x3_Inst201(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6463:6432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst201_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbadbe59),
	.w1(32'hb9f0f76b),
	.w2(32'h39e35838),
	.w3(32'hbb7157c1),
	.w4(32'h3b3aaf81),
	.w5(32'hbbe61409),
	.w6(32'hbb833065),
	.w7(32'h3b27b497),
	.w8(32'hbbdb4892),
)
Conv2D3x3_Inst202(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6495:6464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst202_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3e1008),
	.w1(32'h3b3df1d4),
	.w2(32'h3aa5dd9a),
	.w3(32'hbc2975a8),
	.w4(32'h3939bb34),
	.w5(32'h3b31b21e),
	.w6(32'hbc265be6),
	.w7(32'h3adeca54),
	.w8(32'hba295171),
)
Conv2D3x3_Inst203(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6527:6496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst203_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc25424e),
	.w1(32'hbb837c8d),
	.w2(32'hbb71af5c),
	.w3(32'hbabd8c9a),
	.w4(32'h3b61df71),
	.w5(32'hbb7eb80d),
	.w6(32'hbbc74988),
	.w7(32'h3a822801),
	.w8(32'hbbd0e264),
)
Conv2D3x3_Inst204(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6559:6528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst204_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb10c526),
	.w1(32'hba3da84c),
	.w2(32'h39d9de68),
	.w3(32'hbb30a49b),
	.w4(32'h3a2f89e3),
	.w5(32'hbafb8d97),
	.w6(32'hbb507f04),
	.w7(32'hbabc0139),
	.w8(32'hbb41d634),
)
Conv2D3x3_Inst205(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6591:6560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst205_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3840b9),
	.w1(32'hbb227bac),
	.w2(32'hbbd4177e),
	.w3(32'hbc09edd7),
	.w4(32'h3b8cf358),
	.w5(32'hbb4c9d1e),
	.w6(32'hbc095e33),
	.w7(32'h3ae6c716),
	.w8(32'hbbeccd30),
)
Conv2D3x3_Inst206(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6623:6592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst206_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8a3af5),
	.w1(32'h3b52090b),
	.w2(32'hb9f5974c),
	.w3(32'hbb4712d2),
	.w4(32'h3a842708),
	.w5(32'hbb7af620),
	.w6(32'hbbf397f5),
	.w7(32'hba953a8b),
	.w8(32'hbae7e4f2),
)
Conv2D3x3_Inst207(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6655:6624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst207_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc618217),
	.w1(32'h3b59d7ae),
	.w2(32'hbbb83f54),
	.w3(32'hbbfe4310),
	.w4(32'hbac58adf),
	.w5(32'hbbe5e211),
	.w6(32'h3b044bab),
	.w7(32'hb9576b62),
	.w8(32'hbc1ec986),
)
Conv2D3x3_Inst208(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6687:6656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst208_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9c1fc5a),
	.w1(32'h39998f18),
	.w2(32'h39c896f9),
	.w3(32'hbb48dc53),
	.w4(32'hbaf8cfab),
	.w5(32'hba08a624),
	.w6(32'h3703e2d3),
	.w7(32'hb9fe733f),
	.w8(32'hbadd60ba),
)
Conv2D3x3_Inst209(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6719:6688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst209_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb82216b),
	.w1(32'hbaf7dff4),
	.w2(32'hba9fcba1),
	.w3(32'hbb48a2a8),
	.w4(32'hbb24ef04),
	.w5(32'h3c1ab666),
	.w6(32'hbb15dc74),
	.w7(32'h38bcd29f),
	.w8(32'h3c38e57a),
)
Conv2D3x3_Inst210(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6751:6720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst210_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b17b119),
	.w1(32'h3c100d1f),
	.w2(32'h3bb12c46),
	.w3(32'h3c1b7585),
	.w4(32'h3c1478a6),
	.w5(32'hbb7aedd2),
	.w6(32'h3c03077e),
	.w7(32'h3be20383),
	.w8(32'hbba83e16),
)
Conv2D3x3_Inst211(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6783:6752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst211_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ea150),
	.w1(32'h3ae2ce5a),
	.w2(32'hbbb8bd4d),
	.w3(32'hba91fc53),
	.w4(32'h3ae53060),
	.w5(32'hbc12832e),
	.w6(32'hbb332960),
	.w7(32'h3b4646af),
	.w8(32'hbc27f436),
)
Conv2D3x3_Inst212(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6815:6784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst212_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb833487),
	.w1(32'h3b5ce606),
	.w2(32'hbb42c82d),
	.w3(32'hbb7a3cda),
	.w4(32'h3b9ba21a),
	.w5(32'h3abf30b0),
	.w6(32'hbc7d2efc),
	.w7(32'hbba9f5ed),
	.w8(32'hbbad2cb2),
)
Conv2D3x3_Inst213(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6847:6816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst213_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8bb560),
	.w1(32'hba872f09),
	.w2(32'h3a5c494d),
	.w3(32'hbb9a17d5),
	.w4(32'hbb8a34aa),
	.w5(32'hbb0c2403),
	.w6(32'h3a4eac0e),
	.w7(32'hbb730620),
	.w8(32'hbb31141b),
)
Conv2D3x3_Inst214(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6879:6848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst214_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4396a9),
	.w1(32'hbb7f9d53),
	.w2(32'hbb4c9ed7),
	.w3(32'h3a991b2d),
	.w4(32'h3aed2dad),
	.w5(32'h3a608483),
	.w6(32'hba97ae36),
	.w7(32'hbada9d8d),
	.w8(32'hba1c93a4),
)
Conv2D3x3_Inst215(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6911:6880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst215_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b914bc3),
	.w1(32'hb9eb923b),
	.w2(32'hba766c1c),
	.w3(32'hb9db99af),
	.w4(32'hbb249522),
	.w5(32'h3b29b383),
	.w6(32'hbb0c2187),
	.w7(32'hbb5599db),
	.w8(32'h3b843bb0),
)
Conv2D3x3_Inst216(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6943:6912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst216_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa76e6e),
	.w1(32'h3bff676d),
	.w2(32'hbbd3727d),
	.w3(32'h3bc0f7bc),
	.w4(32'h3b0d7597),
	.w5(32'hbc236d6b),
	.w6(32'h3c5b8618),
	.w7(32'h3b927a5a),
	.w8(32'hbb50ec0e),
)
Conv2D3x3_Inst217(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[6975:6944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst217_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbdb2b44),
	.w1(32'h39982520),
	.w2(32'hbbcb3ee6),
	.w3(32'h3a2bff06),
	.w4(32'hbadc5ec9),
	.w5(32'hbbf845e2),
	.w6(32'h3baefd56),
	.w7(32'hbaf0c459),
	.w8(32'hbc25d127),
)
Conv2D3x3_Inst218(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7007:6976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst218_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc2851c),
	.w1(32'hbb9d3574),
	.w2(32'hbbc12207),
	.w3(32'hbc039ce5),
	.w4(32'hbb61b0bf),
	.w5(32'hbc21c7c2),
	.w6(32'hbb80439d),
	.w7(32'hbafaea18),
	.w8(32'hbc0ee923),
)
Conv2D3x3_Inst219(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7039:7008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst219_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb788cbb),
	.w1(32'h3b2d937c),
	.w2(32'hbb3290ba),
	.w3(32'hbc31ae55),
	.w4(32'h3b1f8b73),
	.w5(32'h3ba1c198),
	.w6(32'hbbf45384),
	.w7(32'hbb47e6c3),
	.w8(32'h3ba773e5),
)
Conv2D3x3_Inst220(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7071:7040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst220_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba580794),
	.w1(32'h3bbfbda4),
	.w2(32'hba97397f),
	.w3(32'hbb483204),
	.w4(32'h3b8b9b75),
	.w5(32'h3a498d67),
	.w6(32'hba7b93a0),
	.w7(32'h3ba52a24),
	.w8(32'hbb8a599e),
)
Conv2D3x3_Inst221(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7103:7072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst221_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb01d009),
	.w1(32'h3bc5a396),
	.w2(32'hbb18ad06),
	.w3(32'h3a6f4def),
	.w4(32'hba90fd34),
	.w5(32'h3b484953),
	.w6(32'h3c240b2b),
	.w7(32'h3a95256d),
	.w8(32'h3b0ce37b),
)
Conv2D3x3_Inst222(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7135:7104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst222_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8bfada),
	.w1(32'h3b324c9b),
	.w2(32'h3a1fd828),
	.w3(32'h3aab3bbb),
	.w4(32'h39168894),
	.w5(32'hbb3a6315),
	.w6(32'h3b80195e),
	.w7(32'hbaf266f9),
	.w8(32'hba0b6ad9),
)
Conv2D3x3_Inst223(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7167:7136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst223_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4c9551),
	.w1(32'hbbeeb116),
	.w2(32'hbabc71c3),
	.w3(32'hbb319b54),
	.w4(32'hbb5a5e4f),
	.w5(32'h3c0b3780),
	.w6(32'hbb624db9),
	.w7(32'h38abba22),
	.w8(32'h3b6ff681),
)
Conv2D3x3_Inst224(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7199:7168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst224_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bd891e2),
	.w1(32'h394040ba),
	.w2(32'hba8ffd4d),
	.w3(32'h3b5b4a63),
	.w4(32'hbab8a0ce),
	.w5(32'h39d63c49),
	.w6(32'h3b372e4d),
	.w7(32'hbaf9e2fa),
	.w8(32'h39735bec),
)
Conv2D3x3_Inst225(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7231:7200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst225_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h384dca92),
	.w1(32'hbaf99d0c),
	.w2(32'hbae8316f),
	.w3(32'hba624451),
	.w4(32'hbb07383a),
	.w5(32'hbac73082),
	.w6(32'hba9e0bb4),
	.w7(32'hbad73dff),
	.w8(32'hba44711a),
)
Conv2D3x3_Inst226(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7263:7232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst226_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5085aa),
	.w1(32'hb93f5765),
	.w2(32'hbb964417),
	.w3(32'h3a45fb1e),
	.w4(32'h3b631f4d),
	.w5(32'hbb01bc61),
	.w6(32'h3a5243f5),
	.w7(32'h3b2e80ca),
	.w8(32'hbb2dedbd),
)
Conv2D3x3_Inst227(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7295:7264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst227_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb623ed0),
	.w1(32'h39eccae4),
	.w2(32'hbaeeb1ce),
	.w3(32'hbb4e0777),
	.w4(32'h3988f06f),
	.w5(32'hbb8ccb40),
	.w6(32'hbb2503f9),
	.w7(32'h399ab315),
	.w8(32'hbb8e03e9),
)
Conv2D3x3_Inst228(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7327:7296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst228_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae748cb),
	.w1(32'hbaa62135),
	.w2(32'hba46cb87),
	.w3(32'hbaa5e5c5),
	.w4(32'hba9690d2),
	.w5(32'h3a4f32d9),
	.w6(32'hba6bb3f3),
	.w7(32'hba678028),
	.w8(32'h3a7c781b),
)
Conv2D3x3_Inst229(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7359:7328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst229_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbab2c515),
	.w1(32'hbb006747),
	.w2(32'hbc0033f0),
	.w3(32'hbb7b095c),
	.w4(32'hbb1abf1d),
	.w5(32'hbbfdc404),
	.w6(32'hbb1e9f74),
	.w7(32'hbab2a59c),
	.w8(32'hbc09fe58),
)
Conv2D3x3_Inst230(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7391:7360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst230_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9eb7d2),
	.w1(32'hba39cac2),
	.w2(32'hbac6782e),
	.w3(32'h3999c0c0),
	.w4(32'hb97bec4a),
	.w5(32'hbb026854),
	.w6(32'hb98c86ef),
	.w7(32'h393bffe2),
	.w8(32'hbb0c5b02),
)
Conv2D3x3_Inst231(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7423:7392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst231_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9a4eb4b),
	.w1(32'hbac87129),
	.w2(32'hbabf8a1c),
	.w3(32'h39382455),
	.w4(32'hb9db4491),
	.w5(32'hb91d8a9d),
	.w6(32'hba827ed8),
	.w7(32'hbaaee902),
	.w8(32'hba7d10a9),
)
Conv2D3x3_Inst232(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7455:7424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst232_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaebc89d),
	.w1(32'h39f3122e),
	.w2(32'hb9d5bdc7),
	.w3(32'hba64688a),
	.w4(32'hb96e570a),
	.w5(32'hbaf78896),
	.w6(32'hba45b078),
	.w7(32'h39d5489f),
	.w8(32'hbae892f6),
)
Conv2D3x3_Inst233(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7487:7456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst233_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb8682749),
	.w1(32'hba712c5b),
	.w2(32'hbab4943f),
	.w3(32'h3a08f5ff),
	.w4(32'h39246e81),
	.w5(32'h3a1b7c17),
	.w6(32'h3a2ca5d1),
	.w7(32'hb9ceb02f),
	.w8(32'h39f8f7d3),
)
Conv2D3x3_Inst234(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7519:7488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst234_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb71e8626),
	.w1(32'hb96ef54a),
	.w2(32'hb8b34b42),
	.w3(32'h3979d054),
	.w4(32'h39d4504d),
	.w5(32'hb839c663),
	.w6(32'hb8a5c8fd),
	.w7(32'hb96365ca),
	.w8(32'hba2550b5),
)
Conv2D3x3_Inst235(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7551:7520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst235_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h39590ee4),
	.w1(32'hba48c433),
	.w2(32'hb929e44f),
	.w3(32'hba8b0859),
	.w4(32'hb9bdf082),
	.w5(32'h38afaac7),
	.w6(32'hbaa2418e),
	.w7(32'hba2ef2b0),
	.w8(32'hba524d37),
)
Conv2D3x3_Inst236(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7583:7552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst236_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb955ecec),
	.w1(32'hba8895e7),
	.w2(32'hba830e3c),
	.w3(32'hba11193a),
	.w4(32'hb9980062),
	.w5(32'h3a117a91),
	.w6(32'hbaed1302),
	.w7(32'hbac9ddfd),
	.w8(32'h3a4c4f92),
)
Conv2D3x3_Inst237(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7615:7584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst237_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb88f59bc),
	.w1(32'h3b3413c6),
	.w2(32'h3a8e522d),
	.w3(32'hbac71bbd),
	.w4(32'h3ad0dd1f),
	.w5(32'hba2097d0),
	.w6(32'hbb0b6be1),
	.w7(32'h39acb39e),
	.w8(32'hbaabf32e),
)
Conv2D3x3_Inst238(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7647:7616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst238_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb173592),
	.w1(32'hbaac27ee),
	.w2(32'hbc2ed1bb),
	.w3(32'hbb04f2c2),
	.w4(32'h37329613),
	.w5(32'hbbc8e7f0),
	.w6(32'hba511006),
	.w7(32'hbabbaa24),
	.w8(32'hbbd22fb3),
)
Conv2D3x3_Inst239(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7679:7648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst239_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae6efb1),
	.w1(32'hba7d2cb6),
	.w2(32'hbb8aaf20),
	.w3(32'h39502c3a),
	.w4(32'h3a5dfdfa),
	.w5(32'hbb44bea9),
	.w6(32'hba90af42),
	.w7(32'h3a68c22b),
	.w8(32'hbb25d35d),
)
Conv2D3x3_Inst240(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7711:7680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst240_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb905d17),
	.w1(32'hbb8070d6),
	.w2(32'hbc010845),
	.w3(32'hbb94e9a9),
	.w4(32'hbb7a5535),
	.w5(32'hbbaf58b9),
	.w6(32'hbb82944b),
	.w7(32'hbb961180),
	.w8(32'hbbcaa31d),
)
Conv2D3x3_Inst241(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7743:7712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst241_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb97ffd80),
	.w1(32'h39c2c44c),
	.w2(32'h3a7e3509),
	.w3(32'h39c79f7b),
	.w4(32'h39124c3f),
	.w5(32'hbb06c4b2),
	.w6(32'h39624ede),
	.w7(32'h39228ba1),
	.w8(32'hbab73ab1),
)
Conv2D3x3_Inst242(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7775:7744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst242_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa42607),
	.w1(32'hbaa3b90f),
	.w2(32'hba937a4f),
	.w3(32'hba9e269a),
	.w4(32'hbaa0b35c),
	.w5(32'h3a91c4a6),
	.w6(32'hbaa0a7de),
	.w7(32'hbac13993),
	.w8(32'h3a6ce101),
)
Conv2D3x3_Inst243(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7807:7776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst243_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a2e88a2),
	.w1(32'h39e52603),
	.w2(32'h3a2af775),
	.w3(32'h3a9932fa),
	.w4(32'h3a9d2c9d),
	.w5(32'hbab14491),
	.w6(32'h3a5ee714),
	.w7(32'h3a8b2790),
	.w8(32'hbac6232f),
)
Conv2D3x3_Inst244(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7839:7808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst244_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba9a2db4),
	.w1(32'hba6e659a),
	.w2(32'hb9c0beed),
	.w3(32'hbaa4e401),
	.w4(32'hba44a91e),
	.w5(32'hb9bd5306),
	.w6(32'hba29324e),
	.w7(32'hb9e38a31),
	.w8(32'hba614e21),
)
Conv2D3x3_Inst245(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7871:7840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst245_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc25d0b),
	.w1(32'hbb828ecf),
	.w2(32'hbbe39620),
	.w3(32'hbb3a23aa),
	.w4(32'hba80a098),
	.w5(32'hbb1448db),
	.w6(32'hbb978870),
	.w7(32'hbb45e3ba),
	.w8(32'hbb718476),
)
Conv2D3x3_Inst246(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7903:7872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst246_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h38d558ed),
	.w1(32'hbabffd06),
	.w2(32'hbaaa8e41),
	.w3(32'hba686d76),
	.w4(32'hba80de69),
	.w5(32'hba98a470),
	.w6(32'hbac791da),
	.w7(32'hbac02803),
	.w8(32'hba294347),
)
Conv2D3x3_Inst247(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7935:7904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst247_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3792d024),
	.w1(32'h3a3e728c),
	.w2(32'hba96c1d9),
	.w3(32'hbace2dca),
	.w4(32'hb98ac5d7),
	.w5(32'h3aa2d12f),
	.w6(32'hba5c551c),
	.w7(32'hba18942a),
	.w8(32'h3a947d8d),
)
Conv2D3x3_Inst248(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7967:7936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst248_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3894d23a),
	.w1(32'hba25de33),
	.w2(32'hb7d98d98),
	.w3(32'hbafb9ee5),
	.w4(32'hb9eb236d),
	.w5(32'hba2a717f),
	.w6(32'hba43eb3e),
	.w7(32'h39ff5dd6),
	.w8(32'hb88c166c),
)
Conv2D3x3_Inst249(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[7999:7968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst249_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h377ea3ff),
	.w1(32'h3acf811b),
	.w2(32'h3b035a4c),
	.w3(32'hba21970f),
	.w4(32'hba8c9f4e),
	.w5(32'h389b623c),
	.w6(32'h392d172e),
	.w7(32'h3921b0a4),
	.w8(32'h39e17f3f),
)
Conv2D3x3_Inst250(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8031:8000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst250_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac0361f),
	.w1(32'hbaadf461),
	.w2(32'hba3847e7),
	.w3(32'hbb0069b5),
	.w4(32'h3a299c6b),
	.w5(32'hba63ac8c),
	.w6(32'hbaf196ac),
	.w7(32'hb990f6cb),
	.w8(32'hbb0a9cd0),
)
Conv2D3x3_Inst251(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8063:8032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst251_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a099c62),
	.w1(32'h3a8c4ed8),
	.w2(32'h3a7ce3b5),
	.w3(32'hb9a31081),
	.w4(32'hb9a214b5),
	.w5(32'h39918365),
	.w6(32'hba7f4dc1),
	.w7(32'hbad83f7f),
	.w8(32'hba5fcd34),
)
Conv2D3x3_Inst252(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8095:8064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst252_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc03adfb),
	.w1(32'hbbaa2279),
	.w2(32'hbc05b124),
	.w3(32'hbb98fc03),
	.w4(32'hbb2a7a3c),
	.w5(32'hba5a2d1d),
	.w6(32'hbb94dc23),
	.w7(32'hbb4237b7),
	.w8(32'hbaad73e8),
)
Conv2D3x3_Inst253(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8127:8096]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst253_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a154436),
	.w1(32'h3994dd6d),
	.w2(32'h3a08d59c),
	.w3(32'h39fce2f7),
	.w4(32'h39f8544e),
	.w5(32'hb6c1d814),
	.w6(32'h39927bc3),
	.w7(32'h39899564),
	.w8(32'hb9d2014e),
)
Conv2D3x3_Inst254(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8159:8128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst254_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaeb6ebc),
	.w1(32'h3ba51f35),
	.w2(32'h3b7730fe),
	.w3(32'hba837bf9),
	.w4(32'h3b21c480),
	.w5(32'h3b496190),
	.w6(32'hbbe4c021),
	.w7(32'hba6310a3),
	.w8(32'h3afec357),
)
Conv2D3x3_Inst255(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[8191:8160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst255_Out),
	.valid_out(valid_out)
);

endmodule