module layer_8_featuremap_195(
	input Clk,
	input Rst,

	input [DATA_WIDTH - 1:0] data_in,
	input valid_in,

	output [DATA_WIDTH - 1:0] data_out,
	output valid_out
);
	parameter DATA_IN_WIDTH = 4096;
	parameter IMG_SIZE = 26;
Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9ca81dc),
	.w1(32'hbc6bc8b2),
	.w2(32'hbc0c8fe8),
	.w3(32'h3a711fe4),
	.w4(32'hbc771bdb),
	.w5(32'hbb92ef00),
	.w6(32'hbc5d2c04),
	.w7(32'hbc49553e),
	.w8(32'hbb23af1b),
)
Conv2D3x3_Inst0(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[31:0]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst0_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0fd486),
	.w1(32'h3c589051),
	.w2(32'h3c49bc6f),
	.w3(32'h3ba9cf3a),
	.w4(32'h3c159f1c),
	.w5(32'h3c1ea78e),
	.w6(32'h3bf6057a),
	.w7(32'h3b9d9ba4),
	.w8(32'h3b751f20),
)
Conv2D3x3_Inst1(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[63:32]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst1_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bf7b8cb),
	.w1(32'h3c21611c),
	.w2(32'h3b7be618),
	.w3(32'h3bd4466e),
	.w4(32'h3c2b14f9),
	.w5(32'h3c58332e),
	.w6(32'h3bb27c2e),
	.w7(32'h39d33b6c),
	.w8(32'h3c2b7362),
)
Conv2D3x3_Inst2(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[95:64]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst2_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b827f7a),
	.w1(32'hbb0a3c51),
	.w2(32'hbb8b1850),
	.w3(32'hbbe75bce),
	.w4(32'hbbddf9f6),
	.w5(32'h3b469d00),
	.w6(32'hb6e68f60),
	.w7(32'hbba1ddda),
	.w8(32'hb9f9141d),
)
Conv2D3x3_Inst3(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[127:96]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst3_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c60b704),
	.w1(32'h3be5eecd),
	.w2(32'h3bfce560),
	.w3(32'hbbaf5158),
	.w4(32'h3b850afa),
	.w5(32'h3b7cbc9f),
	.w6(32'h3a2accac),
	.w7(32'hb97141f7),
	.w8(32'h39d726f7),
)
Conv2D3x3_Inst4(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[159:128]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst4_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aee830f),
	.w1(32'hbc6ec8d4),
	.w2(32'h3d434143),
	.w3(32'h3a2d5922),
	.w4(32'hbc318d03),
	.w5(32'h3d288bdb),
	.w6(32'h3c40496b),
	.w7(32'hbc714a69),
	.w8(32'h3d2991a2),
)
Conv2D3x3_Inst5(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[191:160]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst5_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be93e75),
	.w1(32'hbb5cc176),
	.w2(32'hbbcae4e1),
	.w3(32'hbca7592c),
	.w4(32'hbb1812d4),
	.w5(32'hbb5e2b74),
	.w6(32'h39fa4082),
	.w7(32'hbb3a757c),
	.w8(32'hbb44344d),
)
Conv2D3x3_Inst6(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[223:192]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst6_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be1481b),
	.w1(32'hbc976a9e),
	.w2(32'h3cecb573),
	.w3(32'h3b7f2d18),
	.w4(32'hbc030bba),
	.w5(32'h3d114b58),
	.w6(32'h3c839e6f),
	.w7(32'hbca7c90f),
	.w8(32'h3d083f9c),
)
Conv2D3x3_Inst7(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[255:224]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst7_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c47aa91),
	.w1(32'h3b8eb05b),
	.w2(32'h3bacf698),
	.w3(32'hbc2eb8ed),
	.w4(32'h38cb4886),
	.w5(32'hbb5f05ef),
	.w6(32'hbbc0f62d),
	.w7(32'hbbebd74e),
	.w8(32'hbc19f520),
)
Conv2D3x3_Inst8(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[287:256]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst8_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b80f07e),
	.w1(32'h3be9a4f3),
	.w2(32'hb902b427),
	.w3(32'h3b117d1b),
	.w4(32'h3ba1da30),
	.w5(32'h3c20753d),
	.w6(32'h3c3b324b),
	.w7(32'hba6d9560),
	.w8(32'h3c0b7edc),
)
Conv2D3x3_Inst9(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[319:288]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst9_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb5f2498),
	.w1(32'h3b8b83a1),
	.w2(32'hbc7640a2),
	.w3(32'hbc201247),
	.w4(32'h3b0c1495),
	.w5(32'hbc602afc),
	.w6(32'hbb25e615),
	.w7(32'h3b771e9d),
	.w8(32'hbc08f474),
)
Conv2D3x3_Inst10(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[351:320]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst10_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0dcaf5),
	.w1(32'h3a08f88b),
	.w2(32'hbbca2ab1),
	.w3(32'h39a465c1),
	.w4(32'hb9b4899b),
	.w5(32'h3afa9caf),
	.w6(32'h3a60ebc0),
	.w7(32'hbb1edf28),
	.w8(32'hbb663e2f),
)
Conv2D3x3_Inst11(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[383:352]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst11_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3aa3febd),
	.w1(32'h3c74c71e),
	.w2(32'hbad7c264),
	.w3(32'h3b292575),
	.w4(32'h3b95fac0),
	.w5(32'h3ab08cfb),
	.w6(32'h3b9be519),
	.w7(32'h3c43daf3),
	.w8(32'h3c24df4c),
)
Conv2D3x3_Inst12(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[415:384]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst12_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ac00133),
	.w1(32'hbb8d7965),
	.w2(32'hbb731cb3),
	.w3(32'h39646abd),
	.w4(32'hbc37646e),
	.w5(32'h3c2dc8bb),
	.w6(32'hbb3f1189),
	.w7(32'hbbf48153),
	.w8(32'hb98252a6),
)
Conv2D3x3_Inst13(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[447:416]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst13_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b23f521),
	.w1(32'h3a5c241c),
	.w2(32'hba42e98a),
	.w3(32'hba43cc9e),
	.w4(32'h3aaeec0c),
	.w5(32'hbb2e65c1),
	.w6(32'h3aa01df5),
	.w7(32'hbb18a5e1),
	.w8(32'hbb12a37e),
)
Conv2D3x3_Inst14(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[479:448]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst14_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac387f0),
	.w1(32'hbbd7e74c),
	.w2(32'hbc78aba2),
	.w3(32'hbac61c18),
	.w4(32'h3c325a23),
	.w5(32'hbc674747),
	.w6(32'hbc302d61),
	.w7(32'h3b6a5edb),
	.w8(32'hbc9457ff),
)
Conv2D3x3_Inst15(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[511:480]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst15_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc68ca37),
	.w1(32'h3d02b81b),
	.w2(32'hbc473229),
	.w3(32'h3c715b78),
	.w4(32'hbc21dc48),
	.w5(32'h3ccd9d79),
	.w6(32'h3c03f24b),
	.w7(32'h3ca1f450),
	.w8(32'h3c458811),
)
Conv2D3x3_Inst16(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[543:512]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst16_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d364ba0),
	.w1(32'h3c25aecf),
	.w2(32'hbb4056d6),
	.w3(32'h3c7ea81b),
	.w4(32'h3b862ebb),
	.w5(32'hbb365e3c),
	.w6(32'hbbddf79c),
	.w7(32'h3bb773a7),
	.w8(32'h3a56c25b),
)
Conv2D3x3_Inst17(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[575:544]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst17_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe0174c),
	.w1(32'hbd37e5e0),
	.w2(32'hbb930a7e),
	.w3(32'hbb24d83d),
	.w4(32'hbcb6f2a0),
	.w5(32'hbb37e0cd),
	.w6(32'hbc1f539d),
	.w7(32'hbcb2f3d2),
	.w8(32'hba5ca3a5),
)
Conv2D3x3_Inst18(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[607:576]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst18_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b74f004),
	.w1(32'h3bda3641),
	.w2(32'hbc176a12),
	.w3(32'hbc264644),
	.w4(32'h3aebdd7a),
	.w5(32'hbc6a7dd9),
	.w6(32'h3b8071a5),
	.w7(32'hbbdd5cd5),
	.w8(32'hbc2523dc),
)
Conv2D3x3_Inst19(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[639:608]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst19_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0a5b5e),
	.w1(32'hbbaeb8aa),
	.w2(32'hbc4f0321),
	.w3(32'hbae45b58),
	.w4(32'hb9f3364e),
	.w5(32'hbbe91fae),
	.w6(32'h3ba0fb40),
	.w7(32'hbb250407),
	.w8(32'h3ab5dd87),
)
Conv2D3x3_Inst20(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[671:640]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst20_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae6f144),
	.w1(32'h39d03ae4),
	.w2(32'h3d387288),
	.w3(32'h3bedb313),
	.w4(32'h3cecde03),
	.w5(32'h3c296201),
	.w6(32'hbaa9116a),
	.w7(32'h3c95e767),
	.w8(32'h3c47309e),
)
Conv2D3x3_Inst21(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[703:672]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst21_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc025273),
	.w1(32'h3cb651ab),
	.w2(32'hbcb9fd41),
	.w3(32'h3a287eb4),
	.w4(32'h3c7ee7b1),
	.w5(32'hbd0d85d5),
	.w6(32'hbbfc8506),
	.w7(32'h3c7b9af5),
	.w8(32'hbd32f26c),
)
Conv2D3x3_Inst22(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[735:704]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst22_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa0ee73),
	.w1(32'h3be973e7),
	.w2(32'h3cdb2470),
	.w3(32'h3c7feed1),
	.w4(32'h3c8c4776),
	.w5(32'hbc9453a2),
	.w6(32'hbc63c27e),
	.w7(32'h3c94e148),
	.w8(32'h3b50eb16),
)
Conv2D3x3_Inst23(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[767:736]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst23_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb70d165),
	.w1(32'h3bb708e5),
	.w2(32'h3b83214b),
	.w3(32'h3bcf3fd3),
	.w4(32'h3b97f409),
	.w5(32'h3bac29b7),
	.w6(32'h3aec4d37),
	.w7(32'h3c16a76b),
	.w8(32'h3bb5220a),
)
Conv2D3x3_Inst24(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[799:768]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst24_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ba8be89),
	.w1(32'h3b363853),
	.w2(32'h3c0fcd4f),
	.w3(32'h3ba85ec0),
	.w4(32'h3be62c0d),
	.w5(32'hbc818c7c),
	.w6(32'hbc219a5e),
	.w7(32'hbbc60f9a),
	.w8(32'hbca654df),
)
Conv2D3x3_Inst25(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[831:800]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst25_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc16f231),
	.w1(32'hbc9362b3),
	.w2(32'h3bfbe2de),
	.w3(32'hbb255bc3),
	.w4(32'h39502c44),
	.w5(32'h3a8e15a0),
	.w6(32'h3ab71d44),
	.w7(32'hbbb7bf7e),
	.w8(32'h3c6d2b49),
)
Conv2D3x3_Inst26(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[863:832]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst26_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb3925a),
	.w1(32'hbd160e1d),
	.w2(32'hbdabd9ec),
	.w3(32'hbd31598e),
	.w4(32'hbc984891),
	.w5(32'hbad03b5c),
	.w6(32'hbb044304),
	.w7(32'hbc8043dc),
	.w8(32'hbc9a96bd),
)
Conv2D3x3_Inst27(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[895:864]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst27_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdc884d),
	.w1(32'h3b269885),
	.w2(32'h3b634d6b),
	.w3(32'hbb77226f),
	.w4(32'h3b86af0f),
	.w5(32'h39d33330),
	.w6(32'hbb55d749),
	.w7(32'h3b10352f),
	.w8(32'hbb20817b),
)
Conv2D3x3_Inst28(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[927:896]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst28_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb407aa),
	.w1(32'h3b6d9b36),
	.w2(32'h3bab2943),
	.w3(32'hb83e859c),
	.w4(32'h3bec419e),
	.w5(32'h3c03c5d4),
	.w6(32'h3b215114),
	.w7(32'h3bac6f1c),
	.w8(32'h3c3127a0),
)
Conv2D3x3_Inst29(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[959:928]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst29_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b0a3c8c),
	.w1(32'hb81a0eab),
	.w2(32'hbb8b4e9a),
	.w3(32'h3b8f1b36),
	.w4(32'h38a817a4),
	.w5(32'h3abaa95f),
	.w6(32'h3b4501a9),
	.w7(32'h3bb27648),
	.w8(32'hba69eb2f),
)
Conv2D3x3_Inst30(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[991:960]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst30_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c042b53),
	.w1(32'h3c7ae129),
	.w2(32'h3c0b111b),
	.w3(32'h3ba1d45f),
	.w4(32'h3bc43b0c),
	.w5(32'h3bdc22fe),
	.w6(32'h3b6314cc),
	.w7(32'h3a90160e),
	.w8(32'h3aaf50f4),
)
Conv2D3x3_Inst31(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1023:992]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst31_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3ae30ed4),
	.w1(32'h39c947fb),
	.w2(32'hba7904cd),
	.w3(32'hb9f4a365),
	.w4(32'hbc0caa59),
	.w5(32'hbb2f6745),
	.w6(32'h3af2caa0),
	.w7(32'hbbbf2d99),
	.w8(32'h3b372817),
)
Conv2D3x3_Inst32(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1055:1024]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst32_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c6ee943),
	.w1(32'h3b01d133),
	.w2(32'hbc198d45),
	.w3(32'h3be231b4),
	.w4(32'hbb9252bd),
	.w5(32'hba61444a),
	.w6(32'h3b0257c4),
	.w7(32'hbbaba6c6),
	.w8(32'hbb109eab),
)
Conv2D3x3_Inst33(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1087:1056]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst33_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a9030f6),
	.w1(32'h3c0a300e),
	.w2(32'h3bd10647),
	.w3(32'h3b80be54),
	.w4(32'h3c0cbeac),
	.w5(32'h3b3f5761),
	.w6(32'h3bc962c8),
	.w7(32'h3c062d24),
	.w8(32'h3b35129f),
)
Conv2D3x3_Inst34(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1119:1088]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst34_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb64e56e),
	.w1(32'hbb2ba1b6),
	.w2(32'hbbbcec12),
	.w3(32'hbc042147),
	.w4(32'h37c25e17),
	.w5(32'hbc142732),
	.w6(32'h3b31a5c9),
	.w7(32'hbbed8612),
	.w8(32'h3afb03ad),
)
Conv2D3x3_Inst35(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1151:1120]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst35_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1b02f5),
	.w1(32'h3a430438),
	.w2(32'h3b8126df),
	.w3(32'h3bf6185a),
	.w4(32'hbacd2207),
	.w5(32'hba840755),
	.w6(32'h3b5ffddd),
	.w7(32'h3b22ed5c),
	.w8(32'h3b970b16),
)
Conv2D3x3_Inst36(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1183:1152]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst36_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c247236),
	.w1(32'h3c1b3c1b),
	.w2(32'h3c0e4b46),
	.w3(32'h3bab1a2c),
	.w4(32'h3c24c217),
	.w5(32'h3bbf4f84),
	.w6(32'h3b76a938),
	.w7(32'h3bbd0ffa),
	.w8(32'h3b6dce49),
)
Conv2D3x3_Inst37(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1215:1184]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst37_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba83126d),
	.w1(32'hbc0cc4de),
	.w2(32'h3c844a29),
	.w3(32'h3b07bd17),
	.w4(32'h3bb86a00),
	.w5(32'hbc3987d4),
	.w6(32'hbc744f76),
	.w7(32'h3c54be66),
	.w8(32'hbc876687),
)
Conv2D3x3_Inst38(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1247:1216]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst38_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcab2aa1),
	.w1(32'hbc360cb4),
	.w2(32'hbb88a34e),
	.w3(32'hbc055337),
	.w4(32'hbb6ba275),
	.w5(32'hbc24aa30),
	.w6(32'hbbe00f17),
	.w7(32'hbb89ffc5),
	.w8(32'h3b52c03c),
)
Conv2D3x3_Inst39(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1279:1248]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst39_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc0439c4),
	.w1(32'h3bbc93ca),
	.w2(32'hbafa0435),
	.w3(32'hbc2306ec),
	.w4(32'hbaabe507),
	.w5(32'hbbff4390),
	.w6(32'h3bd5b9ff),
	.w7(32'hbaa203f7),
	.w8(32'hbaa981bb),
)
Conv2D3x3_Inst40(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1311:1280]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst40_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a923ecc),
	.w1(32'h3b78ef3c),
	.w2(32'h39e458b0),
	.w3(32'h3a8987eb),
	.w4(32'h3ae27ec2),
	.w5(32'hba76e848),
	.w6(32'hb888a5b8),
	.w7(32'h3bcbe6f5),
	.w8(32'hbbe9de3b),
)
Conv2D3x3_Inst41(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1343:1312]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst41_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bb5d2e9),
	.w1(32'hb98a66f4),
	.w2(32'h3c0ae16d),
	.w3(32'h3c1a6e7b),
	.w4(32'h3aa11382),
	.w5(32'hbb837ff3),
	.w6(32'hbbc4a8d2),
	.w7(32'hbacd53d2),
	.w8(32'h3937e264),
)
Conv2D3x3_Inst42(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1375:1344]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst42_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b50dbc2),
	.w1(32'hbc9d07ed),
	.w2(32'hbce28628),
	.w3(32'hbb42ab6e),
	.w4(32'hbc300a4b),
	.w5(32'hbc76820b),
	.w6(32'hbc7e8290),
	.w7(32'hbc012810),
	.w8(32'hbc89039d),
)
Conv2D3x3_Inst43(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1407:1376]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst43_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc2fb604),
	.w1(32'hbc14e038),
	.w2(32'hbcbbf74e),
	.w3(32'h3a8aad18),
	.w4(32'hbcbedec7),
	.w5(32'hbc53ebe6),
	.w6(32'h3ab0d40f),
	.w7(32'hbcba6aa3),
	.w8(32'hbb4ca03e),
)
Conv2D3x3_Inst44(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1439:1408]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst44_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c632c83),
	.w1(32'hbb8c7565),
	.w2(32'hbbb8e693),
	.w3(32'h3b077117),
	.w4(32'hbb1f8f26),
	.w5(32'hbb2d33e0),
	.w6(32'hbadd84e5),
	.w7(32'hbbc86510),
	.w8(32'h390a8c5f),
)
Conv2D3x3_Inst45(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1471:1440]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst45_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbac253f4),
	.w1(32'h399e46d3),
	.w2(32'hbc98353b),
	.w3(32'hb9dc930e),
	.w4(32'hba936f77),
	.w5(32'hbc4bea8f),
	.w6(32'hbb832fe9),
	.w7(32'hbc2edb8a),
	.w8(32'hbc4374c9),
)
Conv2D3x3_Inst46(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1503:1472]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst46_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbae6a149),
	.w1(32'hbc4e3894),
	.w2(32'hbb97e69e),
	.w3(32'hbbb616f4),
	.w4(32'h3b9f7921),
	.w5(32'hbc9f26ce),
	.w6(32'hbbb2d3f6),
	.w7(32'hbc394fff),
	.w8(32'h3b398fb2),
)
Conv2D3x3_Inst47(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1535:1504]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst47_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcad5d19),
	.w1(32'hbc5cd721),
	.w2(32'hbc60f7e2),
	.w3(32'hbc35fe73),
	.w4(32'hbb73cd02),
	.w5(32'hbc9110cf),
	.w6(32'hbc809283),
	.w7(32'hbc5504a1),
	.w8(32'h3b4c6c7a),
)
Conv2D3x3_Inst48(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1567:1536]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst48_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbb7353),
	.w1(32'hbba3befb),
	.w2(32'hbc6f796c),
	.w3(32'hbb6f92d8),
	.w4(32'hbb45129e),
	.w5(32'hbba2ee31),
	.w6(32'hba4ec6e7),
	.w7(32'hbc33efd5),
	.w8(32'hbc13e7f3),
)
Conv2D3x3_Inst49(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1599:1568]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst49_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c988adf),
	.w1(32'h3cab5a73),
	.w2(32'h3cc046f2),
	.w3(32'h3cc926b4),
	.w4(32'h3cb4cd25),
	.w5(32'h3cb3d22e),
	.w6(32'h3cb37678),
	.w7(32'h3c9c23a4),
	.w8(32'h3c9337b8),
)
Conv2D3x3_Inst50(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1631:1600]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst50_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8c35b5),
	.w1(32'hbc7b4849),
	.w2(32'hbc634848),
	.w3(32'h3b44d61d),
	.w4(32'hbbfadbd0),
	.w5(32'hbc8dae6c),
	.w6(32'h3b079c54),
	.w7(32'hba9e487a),
	.w8(32'hbc31a8e8),
)
Conv2D3x3_Inst51(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1663:1632]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst51_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bee3e54),
	.w1(32'h3a123f36),
	.w2(32'h3b6c02da),
	.w3(32'h3c136786),
	.w4(32'hbb92396f),
	.w5(32'hbb612991),
	.w6(32'hbbce354b),
	.w7(32'hbc50121f),
	.w8(32'hbc06f869),
)
Conv2D3x3_Inst52(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1695:1664]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst52_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b83ea99),
	.w1(32'hbcc3d803),
	.w2(32'h3cab519d),
	.w3(32'h3b05157a),
	.w4(32'h3a0f7d41),
	.w5(32'hba7c7159),
	.w6(32'hbca0eb15),
	.w7(32'h3ab03ed9),
	.w8(32'hbb7b593b),
)
Conv2D3x3_Inst53(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1727:1696]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst53_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc940b99),
	.w1(32'hbc11eec8),
	.w2(32'hbc2eb5db),
	.w3(32'hbc9d2c3a),
	.w4(32'hbb765abc),
	.w5(32'hba2f27b6),
	.w6(32'h3b4148dc),
	.w7(32'hbbd91dcc),
	.w8(32'hbbd98ee8),
)
Conv2D3x3_Inst54(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1759:1728]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst54_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c0c48e1),
	.w1(32'hba8d5ba7),
	.w2(32'hbc304419),
	.w3(32'h3a6d407b),
	.w4(32'hbb97017b),
	.w5(32'hbad1cbd9),
	.w6(32'h3bd6a56b),
	.w7(32'hbc06c27f),
	.w8(32'hbbb41f9a),
)
Conv2D3x3_Inst55(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1791:1760]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst55_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8c75c6),
	.w1(32'h3cd983a6),
	.w2(32'hbc699490),
	.w3(32'h3c435d8f),
	.w4(32'h3c8d2eb7),
	.w5(32'hbca7bbcb),
	.w6(32'h3baa672a),
	.w7(32'h3cb0bc5c),
	.w8(32'hbc9920c8),
)
Conv2D3x3_Inst56(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1823:1792]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst56_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad0f329),
	.w1(32'hbc15c974),
	.w2(32'hba001add),
	.w3(32'h3c527f30),
	.w4(32'hbb6e091d),
	.w5(32'hbc0a161f),
	.w6(32'hbb3bfb54),
	.w7(32'hba583583),
	.w8(32'hba6087f1),
)
Conv2D3x3_Inst57(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1855:1824]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst57_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b3970ba),
	.w1(32'hbba442a8),
	.w2(32'hbbcb5b18),
	.w3(32'hbb01c87c),
	.w4(32'hbb77564e),
	.w5(32'hbbb63134),
	.w6(32'hbb9d4b0a),
	.w7(32'hbae8841f),
	.w8(32'h388c4508),
)
Conv2D3x3_Inst58(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1887:1856]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst58_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6af283),
	.w1(32'h3c6ac7a9),
	.w2(32'h3d320dbd),
	.w3(32'h39ba3058),
	.w4(32'h3ce431b3),
	.w5(32'hbbcbaf6b),
	.w6(32'hbb00a191),
	.w7(32'h3d1079f7),
	.w8(32'hb7e4039e),
)
Conv2D3x3_Inst59(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1919:1888]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst59_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc831eee),
	.w1(32'hbbf21f61),
	.w2(32'hba5539ef),
	.w3(32'h3c0b0bff),
	.w4(32'hba39dc21),
	.w5(32'hbac3ad5f),
	.w6(32'hbbe435e7),
	.w7(32'hbb354565),
	.w8(32'h3b8deedd),
)
Conv2D3x3_Inst60(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1951:1920]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst60_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3be2a402),
	.w1(32'h3c0709e2),
	.w2(32'hbacd3fd7),
	.w3(32'hbae5d02a),
	.w4(32'h3b88a499),
	.w5(32'h3b2c9dba),
	.w6(32'h3b5b5ee1),
	.w7(32'hb9998053),
	.w8(32'h3b34eb87),
)
Conv2D3x3_Inst61(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[1983:1952]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst61_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c08ff62),
	.w1(32'h3c53550f),
	.w2(32'h3b44fa92),
	.w3(32'h39094bbb),
	.w4(32'hba66ffc9),
	.w5(32'h3c1023b3),
	.w6(32'h3bdc7532),
	.w7(32'hbb1d4890),
	.w8(32'hba09b06b),
)
Conv2D3x3_Inst62(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2015:1984]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst62_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c20069a),
	.w1(32'h3900a430),
	.w2(32'hba2737be),
	.w3(32'h3a0b42d9),
	.w4(32'h3aaf2967),
	.w5(32'hbb9170da),
	.w6(32'h3ab7fa36),
	.w7(32'h3abce3f8),
	.w8(32'h39cca39c),
)
Conv2D3x3_Inst63(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2047:2016]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst63_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaa62af8),
	.w1(32'hb9d48f66),
	.w2(32'hba146b7d),
	.w3(32'hbb701eb3),
	.w4(32'hbb665a2f),
	.w5(32'hbb503b7d),
	.w6(32'hba94470d),
	.w7(32'h3a9362f9),
	.w8(32'hbaa4ed2b),
)
Conv2D3x3_Inst64(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2079:2048]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst64_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b294325),
	.w1(32'hbc5c44d0),
	.w2(32'h3b9d05f8),
	.w3(32'hb90c665a),
	.w4(32'hbb8e1548),
	.w5(32'hbcd50919),
	.w6(32'hbc9b6399),
	.w7(32'hbc125ec2),
	.w8(32'hbb380938),
)
Conv2D3x3_Inst65(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2111:2080]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst65_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba66aac),
	.w1(32'h3bd228ca),
	.w2(32'h3b701d94),
	.w3(32'hbb1e6a85),
	.w4(32'h3b510c44),
	.w5(32'hbb06b63f),
	.w6(32'hbc03acf9),
	.w7(32'h3b835278),
	.w8(32'h3ba8a736),
)
Conv2D3x3_Inst66(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2143:2112]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst66_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8523b0),
	.w1(32'hbb2ac401),
	.w2(32'hbc02bbe6),
	.w3(32'hbbe27d23),
	.w4(32'hbb1cef41),
	.w5(32'hbbf8afd4),
	.w6(32'hbb862b44),
	.w7(32'hbbbe77e0),
	.w8(32'hbb5e6fdc),
)
Conv2D3x3_Inst67(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2175:2144]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst67_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc3d1be0),
	.w1(32'h3c00bff7),
	.w2(32'h3a6ca0b9),
	.w3(32'hba8e9be0),
	.w4(32'hba8e8c25),
	.w5(32'h3c093d8b),
	.w6(32'h3c295c45),
	.w7(32'hbbe1982b),
	.w8(32'h3c229f87),
)
Conv2D3x3_Inst68(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2207:2176]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst68_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cb8cf8f),
	.w1(32'hbb552207),
	.w2(32'hbc0eef9f),
	.w3(32'h3b8b58bc),
	.w4(32'hbbc3a227),
	.w5(32'hbca190b9),
	.w6(32'hbc49a556),
	.w7(32'hbb82cfe8),
	.w8(32'h3a5bed4b),
)
Conv2D3x3_Inst69(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2239:2208]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst69_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc08bbdf),
	.w1(32'hbb0e7e32),
	.w2(32'hbbae0104),
	.w3(32'hbc0f14ef),
	.w4(32'hbab411c0),
	.w5(32'hbb879ffc),
	.w6(32'hbb93b705),
	.w7(32'hbb46855b),
	.w8(32'h3a8585dc),
)
Conv2D3x3_Inst70(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2271:2240]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst70_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bafd712),
	.w1(32'h3baae8dd),
	.w2(32'h3baa0b29),
	.w3(32'h3b8d9e84),
	.w4(32'hbba12637),
	.w5(32'h3c046f87),
	.w6(32'h39b89262),
	.w7(32'hbbe615fe),
	.w8(32'h3b367884),
)
Conv2D3x3_Inst71(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2303:2272]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst71_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c05cb6d),
	.w1(32'h3b255e33),
	.w2(32'hbb037d83),
	.w3(32'hbb40fae6),
	.w4(32'h3b548634),
	.w5(32'h3be7dd4d),
	.w6(32'h398dd7e0),
	.w7(32'hbaeb809f),
	.w8(32'h3c8616b6),
)
Conv2D3x3_Inst72(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2335:2304]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst72_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cbc0f42),
	.w1(32'hbc2dc4fa),
	.w2(32'h3bfd5ff6),
	.w3(32'h3c203839),
	.w4(32'h3b545e5c),
	.w5(32'h3a969926),
	.w6(32'hbbea9482),
	.w7(32'h3937443b),
	.w8(32'h39e03d23),
)
Conv2D3x3_Inst73(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2367:2336]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst73_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbff0444),
	.w1(32'hbb9b918d),
	.w2(32'hbc118519),
	.w3(32'h3ab5e070),
	.w4(32'hbac7a85b),
	.w5(32'hbbee1942),
	.w6(32'hba9b4f0b),
	.w7(32'h3ad532fb),
	.w8(32'hbc487a60),
)
Conv2D3x3_Inst74(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2399:2368]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst74_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbaacb1b0),
	.w1(32'h39db9ed2),
	.w2(32'h3953103d),
	.w3(32'h3c2b3a8f),
	.w4(32'h3c2876cd),
	.w5(32'hbc02590d),
	.w6(32'h38d04311),
	.w7(32'h39a6ce3b),
	.w8(32'hbc866cf8),
)
Conv2D3x3_Inst75(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2431:2400]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst75_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc17fc19),
	.w1(32'hbc011e64),
	.w2(32'hbb847fef),
	.w3(32'hbb8cf98f),
	.w4(32'h3b9c2d82),
	.w5(32'hbc29d181),
	.w6(32'hbc30d72c),
	.w7(32'h3bdd9779),
	.w8(32'hbbed4fcf),
)
Conv2D3x3_Inst76(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2463:2432]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst76_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb4ce047),
	.w1(32'hbbbcedde),
	.w2(32'hbb0eb6b9),
	.w3(32'hba76c03e),
	.w4(32'hba93eadf),
	.w5(32'hbc8211dd),
	.w6(32'hbc09e3a9),
	.w7(32'hbb887d03),
	.w8(32'hbc6bee5f),
)
Conv2D3x3_Inst77(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2495:2464]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst77_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba81f222),
	.w1(32'hbac75e46),
	.w2(32'h39e241fc),
	.w3(32'h3b1ca7da),
	.w4(32'hba4844ba),
	.w5(32'hbb498003),
	.w6(32'hbb51de50),
	.w7(32'hbb851247),
	.w8(32'h3ab4918a),
)
Conv2D3x3_Inst78(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2527:2496]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst78_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bbbc80d),
	.w1(32'hbc2562fb),
	.w2(32'hbca072c5),
	.w3(32'h3b48ac8b),
	.w4(32'hbc39481e),
	.w5(32'h3b74e444),
	.w6(32'hbb44f157),
	.w7(32'hbc87798d),
	.w8(32'h3c1e30a7),
)
Conv2D3x3_Inst79(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2559:2528]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst79_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3fd815),
	.w1(32'h3ae708a6),
	.w2(32'hbabafba3),
	.w3(32'h3b612dea),
	.w4(32'hbc0f6b70),
	.w5(32'h3b079718),
	.w6(32'h3b47d9aa),
	.w7(32'hbba3d6e6),
	.w8(32'h3b854b65),
)
Conv2D3x3_Inst80(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2591:2560]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst80_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a77bb8c),
	.w1(32'h3ba9a72d),
	.w2(32'h3b8a923e),
	.w3(32'hbbc5f844),
	.w4(32'hbaee4b92),
	.w5(32'h3bca5978),
	.w6(32'hb9f86044),
	.w7(32'hbc487126),
	.w8(32'h39dc124f),
)
Conv2D3x3_Inst81(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2623:2592]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst81_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b81b956),
	.w1(32'hbba83bdf),
	.w2(32'h3c34a796),
	.w3(32'hb9ef5785),
	.w4(32'h3b0b2a3c),
	.w5(32'hbc26acb7),
	.w6(32'hbc45d247),
	.w7(32'h3be0353e),
	.w8(32'hbbcb531e),
)
Conv2D3x3_Inst82(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2655:2624]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst82_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb61ace),
	.w1(32'hbc3329f7),
	.w2(32'h3d1a15b9),
	.w3(32'h3c0e2b3a),
	.w4(32'hbb7b80e4),
	.w5(32'h3d2d02bb),
	.w6(32'h3c897d60),
	.w7(32'h3b32a32f),
	.w8(32'h3d0adf8b),
)
Conv2D3x3_Inst83(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2687:2656]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst83_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c3b9f85),
	.w1(32'h3c0eaca0),
	.w2(32'hbbad21bf),
	.w3(32'hbc02cdc2),
	.w4(32'hbbd7f4b7),
	.w5(32'h3a063c6f),
	.w6(32'hba8cb7a1),
	.w7(32'hbca1e5ad),
	.w8(32'hbc07337f),
)
Conv2D3x3_Inst84(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2719:2688]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst84_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cae7e1c),
	.w1(32'hbbbf9969),
	.w2(32'h3a960325),
	.w3(32'h3bc6d7d4),
	.w4(32'h3b80e239),
	.w5(32'hbb8a2e27),
	.w6(32'hbabceb23),
	.w7(32'hbc446d74),
	.w8(32'h3bc80599),
)
Conv2D3x3_Inst85(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2751:2720]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst85_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c273737),
	.w1(32'h3915828d),
	.w2(32'h3b5508e1),
	.w3(32'h3bc2907f),
	.w4(32'h3a252e0b),
	.w5(32'h3b900799),
	.w6(32'hbabc637c),
	.w7(32'h3a66c7f6),
	.w8(32'h3a07a235),
)
Conv2D3x3_Inst86(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2783:2752]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst86_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3aaa83),
	.w1(32'h3b208b12),
	.w2(32'hba7ec45b),
	.w3(32'hbb30ad7d),
	.w4(32'hbabbfc9d),
	.w5(32'h3abc0370),
	.w6(32'h3b4af828),
	.w7(32'h3b9e6e6a),
	.w8(32'hba93ccc7),
)
Conv2D3x3_Inst87(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2815:2784]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst87_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b88e5e6),
	.w1(32'h3a9f3255),
	.w2(32'h3aa10c79),
	.w3(32'h3b2ee2fc),
	.w4(32'h3b60d7b6),
	.w5(32'h3baa9e9b),
	.w6(32'h3ae56cc6),
	.w7(32'h3a8df484),
	.w8(32'h3ad68b19),
)
Conv2D3x3_Inst88(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2847:2816]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst88_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bccd99a),
	.w1(32'hbb9f2749),
	.w2(32'h3b33e8ff),
	.w3(32'h3bb0e3f9),
	.w4(32'hbb4b934e),
	.w5(32'hbc00b883),
	.w6(32'hbb86ea41),
	.w7(32'h3b034166),
	.w8(32'hbaaa3bb3),
)
Conv2D3x3_Inst89(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2879:2848]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst89_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc223396),
	.w1(32'h3ba4d23a),
	.w2(32'hb9c02f3c),
	.w3(32'hba83ed3f),
	.w4(32'hbac8e08c),
	.w5(32'h3c35d700),
	.w6(32'h3c17acf2),
	.w7(32'h3b230b95),
	.w8(32'h3c172782),
)
Conv2D3x3_Inst90(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2911:2880]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst90_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c582ded),
	.w1(32'hb9c55f71),
	.w2(32'hbc19a259),
	.w3(32'hbbfd3200),
	.w4(32'h391ba207),
	.w5(32'hb90de0ad),
	.w6(32'hbc0702b8),
	.w7(32'hbb4352c7),
	.w8(32'hbc1ac9c9),
)
Conv2D3x3_Inst91(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2943:2912]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst91_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbe975db),
	.w1(32'h3b102a2b),
	.w2(32'h3b6c5e35),
	.w3(32'hb9504448),
	.w4(32'hbaeddfb7),
	.w5(32'hb90c3643),
	.w6(32'h3a8fd40d),
	.w7(32'h3aca875d),
	.w8(32'hb857552c),
)
Conv2D3x3_Inst92(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[2975:2944]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst92_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b2ef825),
	.w1(32'hbbb89763),
	.w2(32'hbba11b95),
	.w3(32'hbb20ec6d),
	.w4(32'hbbed3b2e),
	.w5(32'hbbdbf087),
	.w6(32'hbc0a5b85),
	.w7(32'hbc130dbb),
	.w8(32'hbc2c09ee),
)
Conv2D3x3_Inst93(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3007:2976]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst93_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb1c6e53),
	.w1(32'hbc78f390),
	.w2(32'h3c5f6f91),
	.w3(32'hbb4e3005),
	.w4(32'hbbb99f9d),
	.w5(32'h3c8793c8),
	.w6(32'h3a73c76d),
	.w7(32'hbbd5bcbd),
	.w8(32'h3c8fbb5c),
)
Conv2D3x3_Inst94(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3039:3008]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst94_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba4e3d6f),
	.w1(32'hbc178a9f),
	.w2(32'hbbff8567),
	.w3(32'hbc718c94),
	.w4(32'hbb61c08b),
	.w5(32'hbb357c49),
	.w6(32'hbb85b61b),
	.w7(32'hbbc1ab0a),
	.w8(32'hbb38607c),
)
Conv2D3x3_Inst95(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3071:3040]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst95_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c693688),
	.w1(32'hba2bd503),
	.w2(32'h3c1a7f5d),
	.w3(32'h3c4af33d),
	.w4(32'h3c3e2dd3),
	.w5(32'hbc838684),
	.w6(32'hbc11dae4),
	.w7(32'h3c571e0d),
	.w8(32'hbcab5a11),
)
Conv2D3x3_Inst96(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3103:3072]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst96_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcbc5bdc),
	.w1(32'hbc546991),
	.w2(32'h3c8f9d34),
	.w3(32'hbc751418),
	.w4(32'h3c473c9f),
	.w5(32'hbbfe0a6a),
	.w6(32'hbce0e09e),
	.w7(32'h3c09eee4),
	.w8(32'hbc9f23df),
)
Conv2D3x3_Inst97(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3135:3104]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst97_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcf1a092),
	.w1(32'hbb8de9dd),
	.w2(32'hbbde6e48),
	.w3(32'hbc642d1a),
	.w4(32'h3ba5e06e),
	.w5(32'hbc6d2dcd),
	.w6(32'hbc2ecadc),
	.w7(32'h3b9c8c8e),
	.w8(32'hbca803d6),
)
Conv2D3x3_Inst98(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3167:3136]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst98_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbc8a3e23),
	.w1(32'hbbcfa737),
	.w2(32'hbb82fc36),
	.w3(32'hbb95a1a0),
	.w4(32'hbbef750c),
	.w5(32'h3c1474c5),
	.w6(32'hbc263c22),
	.w7(32'h3bab82f8),
	.w8(32'hbb881acf),
)
Conv2D3x3_Inst99(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3199:3168]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst99_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb7b605e),
	.w1(32'hbb9a81f1),
	.w2(32'hbc0cf29f),
	.w3(32'hbc3507e2),
	.w4(32'hbc3aed8e),
	.w5(32'hbca51926),
	.w6(32'hbbc1ca06),
	.w7(32'h3b4ac276),
	.w8(32'hbb3c992f),
)
Conv2D3x3_Inst100(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3231:3200]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst100_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb9c8c74),
	.w1(32'hba7b03f4),
	.w2(32'hbc8d9176),
	.w3(32'h3be77f00),
	.w4(32'hbced8097),
	.w5(32'h3cfc771d),
	.w6(32'h3cf6768b),
	.w7(32'hbd1d5684),
	.w8(32'hbadbc505),
)
Conv2D3x3_Inst101(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3263:3232]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst101_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3d05a6d8),
	.w1(32'hbb3ce54f),
	.w2(32'h3ad3e420),
	.w3(32'hbb88b803),
	.w4(32'hbbac2372),
	.w5(32'hba8f6ec6),
	.w6(32'hb9e9b0fa),
	.w7(32'hbb97b1c8),
	.w8(32'hbc0e87e1),
)
Conv2D3x3_Inst102(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3295:3264]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst102_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb8ace13),
	.w1(32'h3cee407e),
	.w2(32'hbbd60447),
	.w3(32'hbb884196),
	.w4(32'h3c4572d3),
	.w5(32'hbc7543b8),
	.w6(32'hbc0d03e2),
	.w7(32'h3cfddc4b),
	.w8(32'hbc246740),
)
Conv2D3x3_Inst103(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3327:3296]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst103_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bdf3ba3),
	.w1(32'h3d1388a4),
	.w2(32'hbb422dc2),
	.w3(32'h3c510ca9),
	.w4(32'h3ccc937e),
	.w5(32'h3c7459c3),
	.w6(32'h3c35dbcf),
	.w7(32'h3c9c78e0),
	.w8(32'hbb72c8b6),
)
Conv2D3x3_Inst104(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3359:3328]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst104_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3cc914af),
	.w1(32'hbbb7ed63),
	.w2(32'hbc18584f),
	.w3(32'h3cb141f8),
	.w4(32'hbc21d29c),
	.w5(32'hbc41cc3f),
	.w6(32'hbc5e34ab),
	.w7(32'hbc56031b),
	.w8(32'hbc0c7916),
)
Conv2D3x3_Inst105(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3391:3360]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst105_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a8bc7ed),
	.w1(32'hbb79ec88),
	.w2(32'hbbde112f),
	.w3(32'hb9b25814),
	.w4(32'hbb10b883),
	.w5(32'hbc409a98),
	.w6(32'hbbc23ef8),
	.w7(32'hbc1c55df),
	.w8(32'hbc88cb52),
)
Conv2D3x3_Inst106(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3423:3392]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst106_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbb92264),
	.w1(32'hb961bf92),
	.w2(32'hba3b8a66),
	.w3(32'hbb9a7bf2),
	.w4(32'hbaf4d5c8),
	.w5(32'hbb94027f),
	.w6(32'hbb9ce9b8),
	.w7(32'hbc345d2c),
	.w8(32'hba5cb4ce),
)
Conv2D3x3_Inst107(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3455:3424]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst107_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb98db03f),
	.w1(32'h3b934ae0),
	.w2(32'h3b743d90),
	.w3(32'h3a7e499a),
	.w4(32'h3bd1abe5),
	.w5(32'h3c09112b),
	.w6(32'h3bcedd29),
	.w7(32'h3b95e5de),
	.w8(32'h3b34c803),
)
Conv2D3x3_Inst108(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3487:3456]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst108_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c1e5694),
	.w1(32'h3bc5872d),
	.w2(32'h3bbd8e0c),
	.w3(32'h3c05957f),
	.w4(32'h3ad338cf),
	.w5(32'h3af720f2),
	.w6(32'h39fd70f5),
	.w7(32'h398148cc),
	.w8(32'hbad7d03a),
)
Conv2D3x3_Inst109(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3519:3488]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst109_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hb9b7e391),
	.w1(32'h3bbb7b1a),
	.w2(32'h3b7a46fa),
	.w3(32'hbb56a406),
	.w4(32'h3b868018),
	.w5(32'h3c1593ea),
	.w6(32'h395fc355),
	.w7(32'h3b1f777b),
	.w8(32'hba12c9ac),
)
Conv2D3x3_Inst110(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3551:3520]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst110_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba3d97de),
	.w1(32'h3b852190),
	.w2(32'h3be10e30),
	.w3(32'hbb528ee7),
	.w4(32'h3b9c953e),
	.w5(32'h3b986065),
	.w6(32'h3b3eeaa8),
	.w7(32'h3be7e348),
	.w8(32'h3bebb6b3),
)
Conv2D3x3_Inst111(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3583:3552]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst111_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3bcf5ea1),
	.w1(32'h3c148742),
	.w2(32'hb776d78b),
	.w3(32'h3bba157e),
	.w4(32'h3c12c9b7),
	.w5(32'h3ad78184),
	.w6(32'h3bb3f831),
	.w7(32'h3c5363b6),
	.w8(32'h3c542d84),
)
Conv2D3x3_Inst112(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3615:3584]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst112_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbba74f51),
	.w1(32'h3be183e2),
	.w2(32'hbaee589e),
	.w3(32'hba8162dc),
	.w4(32'hbbc1a991),
	.w5(32'hba29f93c),
	.w6(32'hbb4be2cc),
	.w7(32'h3b9dec30),
	.w8(32'h3bdbf1a4),
)
Conv2D3x3_Inst113(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3647:3616]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst113_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbc7612a),
	.w1(32'hbb4648f5),
	.w2(32'h3aac87b3),
	.w3(32'hbae8929a),
	.w4(32'h3b6b36d3),
	.w5(32'h39810da6),
	.w6(32'hbb648b45),
	.w7(32'hbb117cae),
	.w8(32'h3b86d397),
)
Conv2D3x3_Inst114(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3679:3648]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst114_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b8b3353),
	.w1(32'hba7a2c86),
	.w2(32'h3a30557c),
	.w3(32'h3aafa744),
	.w4(32'hbb54f2d4),
	.w5(32'h390bfa86),
	.w6(32'hba4fe7c0),
	.w7(32'hba468b69),
	.w8(32'hbacdc602),
)
Conv2D3x3_Inst115(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3711:3680]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst115_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hba8af071),
	.w1(32'hbb463956),
	.w2(32'hba79d670),
	.w3(32'hbb217827),
	.w4(32'h3ad7491e),
	.w5(32'hba2fd0a2),
	.w6(32'h3a65990d),
	.w7(32'h3aa9fa62),
	.w8(32'h3b8174b5),
)
Conv2D3x3_Inst116(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3743:3712]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst116_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b6db6ea),
	.w1(32'h3bdba2af),
	.w2(32'hbb44810d),
	.w3(32'h3b93eecc),
	.w4(32'h3ae9b433),
	.w5(32'h3bf40c9f),
	.w6(32'h3b2131db),
	.w7(32'hbaa73cd0),
	.w8(32'h3ba4097d),
)
Conv2D3x3_Inst117(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3775:3744]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst117_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b4e3fc7),
	.w1(32'hbb3389ed),
	.w2(32'h3748c2d4),
	.w3(32'h3a39bb25),
	.w4(32'hbb9d2a54),
	.w5(32'h3b6232e6),
	.w6(32'h3bd700e7),
	.w7(32'hbc6a05a1),
	.w8(32'h3aa4eadd),
)
Conv2D3x3_Inst118(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3807:3776]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst118_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b84fea2),
	.w1(32'hb98d1587),
	.w2(32'hbb4675c3),
	.w3(32'hbb254726),
	.w4(32'h3b841d5b),
	.w5(32'hbc260998),
	.w6(32'h38417cfd),
	.w7(32'h3b7a7265),
	.w8(32'hbc169361),
)
Conv2D3x3_Inst119(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3839:3808]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst119_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbbd28166),
	.w1(32'h3beb4795),
	.w2(32'h39e18629),
	.w3(32'h3c294521),
	.w4(32'h3bd136df),
	.w5(32'h3c960862),
	.w6(32'h3cc0819c),
	.w7(32'hba8fcfb2),
	.w8(32'h3bd588cf),
)
Conv2D3x3_Inst120(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3871:3840]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst120_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3b51e0da),
	.w1(32'hbbc39584),
	.w2(32'hbc87bd87),
	.w3(32'h3c11b5f6),
	.w4(32'hbb9d8671),
	.w5(32'hbc155423),
	.w6(32'h3b9273ba),
	.w7(32'hbbe3b712),
	.w8(32'hb9a83c88),
)
Conv2D3x3_Inst121(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3903:3872]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst121_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb3cfbaf),
	.w1(32'hbb272afe),
	.w2(32'h39d430f3),
	.w3(32'hbc095d6f),
	.w4(32'hbade2aec),
	.w5(32'h3b2e2917),
	.w6(32'hbb3aae81),
	.w7(32'hba816d17),
	.w8(32'h39da59b2),
)
Conv2D3x3_Inst122(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3935:3904]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst122_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbb277cbb),
	.w1(32'h3c16d3c9),
	.w2(32'h3b5e7e14),
	.w3(32'hbb2ca150),
	.w4(32'h3bd0eea7),
	.w5(32'h3aa5d05c),
	.w6(32'h3a41ce03),
	.w7(32'h3c36a20f),
	.w8(32'h3bea4aa5),
)
Conv2D3x3_Inst123(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3967:3936]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst123_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3a58cd53),
	.w1(32'h3bb036bf),
	.w2(32'h3c47e920),
	.w3(32'h3aebd3ff),
	.w4(32'hba600b26),
	.w5(32'h3c85f652),
	.w6(32'h3c8b58b7),
	.w7(32'h3b782253),
	.w8(32'h3c7e222c),
)
Conv2D3x3_Inst124(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[3999:3968]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst124_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'h3c8ca4c6),
	.w1(32'h3ad4b040),
	.w2(32'h39d8bf9f),
	.w3(32'hbbee5827),
	.w4(32'h3b3c1639),
	.w5(32'hbcae72fb),
	.w6(32'hbc5dc36e),
	.w7(32'hbaeca9a8),
	.w8(32'h3c0051ee),
)
Conv2D3x3_Inst125(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4031:4000]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst125_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbcd7a675),
	.w1(32'h3b04f095),
	.w2(32'h3a868041),
	.w3(32'hbb1e5ea7),
	.w4(32'h3b56c472),
	.w5(32'hbab2e22b),
	.w6(32'h3bd88857),
	.w7(32'hba46cf07),
	.w8(32'h3b42ad38),
)
Conv2D3x3_Inst126(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4063:4032]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst126_Out),
	.valid_out(valid_out)
);

Conv2D3x3 #(
	.IMG_SIZE(IMG_SIZE)
	.w0(32'hbad5ae2d),
	.w1(32'h3a91765c),
	.w2(32'h3b93fe2b),
	.w3(32'hbb3ef10a),
	.w4(32'h3aff8302),
	.w5(32'hbb3debb1),
	.w6(32'hbbec0f70),
	.w7(32'hbc5715f9),
	.w8(32'hbbdcc8c3),
)
Conv2D3x3_Inst127(
	.Clk(Clk),
	.Rst(Rst),
	.data_in(data_in[4095:4064]),
	.valid_in(valid_in),
	.data_out(Conv2D3x3_Inst127_Out),
	.valid_out(valid_out)
);

endmodule